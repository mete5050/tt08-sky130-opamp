magic
tech sky130B
magscale 1 2
timestamp 1768735973
<< nwell >>
rect -710 -664 710 698
<< pmos >>
rect -616 -564 -416 636
rect -358 -564 -158 636
rect -100 -564 100 636
rect 158 -564 358 636
rect 416 -564 616 636
<< pdiff >>
rect -674 624 -616 636
rect -674 -552 -662 624
rect -628 -552 -616 624
rect -674 -564 -616 -552
rect -416 624 -358 636
rect -416 -552 -404 624
rect -370 -552 -358 624
rect -416 -564 -358 -552
rect -158 624 -100 636
rect -158 -552 -146 624
rect -112 -552 -100 624
rect -158 -564 -100 -552
rect 100 624 158 636
rect 100 -552 112 624
rect 146 -552 158 624
rect 100 -564 158 -552
rect 358 624 416 636
rect 358 -552 370 624
rect 404 -552 416 624
rect 358 -564 416 -552
rect 616 624 674 636
rect 616 -552 628 624
rect 662 -552 674 624
rect 616 -564 674 -552
<< pdiffc >>
rect -662 -552 -628 624
rect -404 -552 -370 624
rect -146 -552 -112 624
rect 112 -552 146 624
rect 370 -552 404 624
rect 628 -552 662 624
<< poly >>
rect -616 636 -416 662
rect -358 636 -158 662
rect -100 636 100 662
rect 158 636 358 662
rect 416 636 616 662
rect -616 -611 -416 -564
rect -616 -645 -600 -611
rect -432 -645 -416 -611
rect -616 -661 -416 -645
rect -358 -611 -158 -564
rect -358 -645 -342 -611
rect -174 -645 -158 -611
rect -358 -661 -158 -645
rect -100 -611 100 -564
rect -100 -645 -84 -611
rect 84 -645 100 -611
rect -100 -661 100 -645
rect 158 -611 358 -564
rect 158 -645 174 -611
rect 342 -645 358 -611
rect 158 -661 358 -645
rect 416 -611 616 -564
rect 416 -645 432 -611
rect 600 -645 616 -611
rect 416 -661 616 -645
<< polycont >>
rect -600 -645 -432 -611
rect -342 -645 -174 -611
rect -84 -645 84 -611
rect 174 -645 342 -611
rect 432 -645 600 -611
<< locali >>
rect -662 624 -628 640
rect -662 -568 -628 -552
rect -404 624 -370 640
rect -404 -568 -370 -552
rect -146 624 -112 640
rect -146 -568 -112 -552
rect 112 624 146 640
rect 112 -568 146 -552
rect 370 624 404 640
rect 370 -568 404 -552
rect 628 624 662 640
rect 628 -568 662 -552
rect -616 -645 -600 -611
rect -432 -645 -416 -611
rect -358 -645 -342 -611
rect -174 -645 -158 -611
rect -100 -645 -84 -611
rect 84 -645 100 -611
rect 158 -645 174 -611
rect 342 -645 358 -611
rect 416 -645 432 -611
rect 600 -645 616 -611
<< viali >>
rect -662 -552 -628 624
rect -404 -552 -370 624
rect -146 -552 -112 624
rect 112 -552 146 624
rect 370 -552 404 624
rect 628 -552 662 624
rect -600 -645 -432 -611
rect -342 -645 -174 -611
rect -84 -645 84 -611
rect 174 -645 342 -611
rect 432 -645 600 -611
<< metal1 >>
rect -668 624 -622 636
rect -668 -552 -662 624
rect -628 -552 -622 624
rect -668 -564 -622 -552
rect -410 624 -364 636
rect -410 -552 -404 624
rect -370 -552 -364 624
rect -410 -564 -364 -552
rect -152 624 -106 636
rect -152 -552 -146 624
rect -112 -552 -106 624
rect -152 -564 -106 -552
rect 106 624 152 636
rect 106 -552 112 624
rect 146 -552 152 624
rect 106 -564 152 -552
rect 364 624 410 636
rect 364 -552 370 624
rect 404 -552 410 624
rect 364 -564 410 -552
rect 622 624 668 636
rect 622 -552 628 624
rect 662 -552 668 624
rect 622 -564 668 -552
rect -612 -611 -420 -605
rect -612 -645 -600 -611
rect -432 -645 -420 -611
rect -612 -651 -420 -645
rect -354 -611 -162 -605
rect -354 -645 -342 -611
rect -174 -645 -162 -611
rect -354 -651 -162 -645
rect -96 -611 96 -605
rect -96 -645 -84 -611
rect 84 -645 96 -611
rect -96 -651 96 -645
rect 162 -611 354 -605
rect 162 -645 174 -611
rect 342 -645 354 -611
rect 162 -651 354 -645
rect 420 -611 612 -605
rect 420 -645 432 -611
rect 600 -645 612 -611
rect 420 -651 612 -645
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
