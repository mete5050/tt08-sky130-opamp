magic
tech sky130B
magscale 1 2
timestamp 1768734963
<< nwell >>
rect -1457 -819 1457 819
<< pmos >>
rect -1261 -600 -1061 600
rect -1003 -600 -803 600
rect -745 -600 -545 600
rect -487 -600 -287 600
rect -229 -600 -29 600
rect 29 -600 229 600
rect 287 -600 487 600
rect 545 -600 745 600
rect 803 -600 1003 600
rect 1061 -600 1261 600
<< pdiff >>
rect -1319 588 -1261 600
rect -1319 -588 -1307 588
rect -1273 -588 -1261 588
rect -1319 -600 -1261 -588
rect -1061 588 -1003 600
rect -1061 -588 -1049 588
rect -1015 -588 -1003 588
rect -1061 -600 -1003 -588
rect -803 588 -745 600
rect -803 -588 -791 588
rect -757 -588 -745 588
rect -803 -600 -745 -588
rect -545 588 -487 600
rect -545 -588 -533 588
rect -499 -588 -487 588
rect -545 -600 -487 -588
rect -287 588 -229 600
rect -287 -588 -275 588
rect -241 -588 -229 588
rect -287 -600 -229 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 229 588 287 600
rect 229 -588 241 588
rect 275 -588 287 588
rect 229 -600 287 -588
rect 487 588 545 600
rect 487 -588 499 588
rect 533 -588 545 588
rect 487 -600 545 -588
rect 745 588 803 600
rect 745 -588 757 588
rect 791 -588 803 588
rect 745 -600 803 -588
rect 1003 588 1061 600
rect 1003 -588 1015 588
rect 1049 -588 1061 588
rect 1003 -600 1061 -588
rect 1261 588 1319 600
rect 1261 -588 1273 588
rect 1307 -588 1319 588
rect 1261 -600 1319 -588
<< pdiffc >>
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
<< nsubdiff >>
rect -1421 749 -1325 783
rect 1325 749 1421 783
rect -1421 687 -1387 749
rect 1387 687 1421 749
rect -1421 -749 -1387 -687
rect 1387 -749 1421 -687
rect -1421 -783 -1325 -749
rect 1325 -783 1421 -749
<< nsubdiffcont >>
rect -1325 749 1325 783
rect -1421 -687 -1387 687
rect 1387 -687 1421 687
rect -1325 -783 1325 -749
<< poly >>
rect -1261 681 -1061 697
rect -1261 647 -1245 681
rect -1077 647 -1061 681
rect -1261 600 -1061 647
rect -1003 681 -803 697
rect -1003 647 -987 681
rect -819 647 -803 681
rect -1003 600 -803 647
rect -745 681 -545 697
rect -745 647 -729 681
rect -561 647 -545 681
rect -745 600 -545 647
rect -487 681 -287 697
rect -487 647 -471 681
rect -303 647 -287 681
rect -487 600 -287 647
rect -229 681 -29 697
rect -229 647 -213 681
rect -45 647 -29 681
rect -229 600 -29 647
rect 29 681 229 697
rect 29 647 45 681
rect 213 647 229 681
rect 29 600 229 647
rect 287 681 487 697
rect 287 647 303 681
rect 471 647 487 681
rect 287 600 487 647
rect 545 681 745 697
rect 545 647 561 681
rect 729 647 745 681
rect 545 600 745 647
rect 803 681 1003 697
rect 803 647 819 681
rect 987 647 1003 681
rect 803 600 1003 647
rect 1061 681 1261 697
rect 1061 647 1077 681
rect 1245 647 1261 681
rect 1061 600 1261 647
rect -1261 -647 -1061 -600
rect -1261 -681 -1245 -647
rect -1077 -681 -1061 -647
rect -1261 -697 -1061 -681
rect -1003 -647 -803 -600
rect -1003 -681 -987 -647
rect -819 -681 -803 -647
rect -1003 -697 -803 -681
rect -745 -647 -545 -600
rect -745 -681 -729 -647
rect -561 -681 -545 -647
rect -745 -697 -545 -681
rect -487 -647 -287 -600
rect -487 -681 -471 -647
rect -303 -681 -287 -647
rect -487 -697 -287 -681
rect -229 -647 -29 -600
rect -229 -681 -213 -647
rect -45 -681 -29 -647
rect -229 -697 -29 -681
rect 29 -647 229 -600
rect 29 -681 45 -647
rect 213 -681 229 -647
rect 29 -697 229 -681
rect 287 -647 487 -600
rect 287 -681 303 -647
rect 471 -681 487 -647
rect 287 -697 487 -681
rect 545 -647 745 -600
rect 545 -681 561 -647
rect 729 -681 745 -647
rect 545 -697 745 -681
rect 803 -647 1003 -600
rect 803 -681 819 -647
rect 987 -681 1003 -647
rect 803 -697 1003 -681
rect 1061 -647 1261 -600
rect 1061 -681 1077 -647
rect 1245 -681 1261 -647
rect 1061 -697 1261 -681
<< polycont >>
rect -1245 647 -1077 681
rect -987 647 -819 681
rect -729 647 -561 681
rect -471 647 -303 681
rect -213 647 -45 681
rect 45 647 213 681
rect 303 647 471 681
rect 561 647 729 681
rect 819 647 987 681
rect 1077 647 1245 681
rect -1245 -681 -1077 -647
rect -987 -681 -819 -647
rect -729 -681 -561 -647
rect -471 -681 -303 -647
rect -213 -681 -45 -647
rect 45 -681 213 -647
rect 303 -681 471 -647
rect 561 -681 729 -647
rect 819 -681 987 -647
rect 1077 -681 1245 -647
<< locali >>
rect -1421 749 -1325 783
rect 1325 749 1421 783
rect -1421 687 -1387 749
rect 1387 687 1421 749
rect -1261 647 -1245 681
rect -1077 647 -1061 681
rect -1003 647 -987 681
rect -819 647 -803 681
rect -745 647 -729 681
rect -561 647 -545 681
rect -487 647 -471 681
rect -303 647 -287 681
rect -229 647 -213 681
rect -45 647 -29 681
rect 29 647 45 681
rect 213 647 229 681
rect 287 647 303 681
rect 471 647 487 681
rect 545 647 561 681
rect 729 647 745 681
rect 803 647 819 681
rect 987 647 1003 681
rect 1061 647 1077 681
rect 1245 647 1261 681
rect -1307 588 -1273 604
rect -1307 -604 -1273 -588
rect -1049 588 -1015 604
rect -1049 -604 -1015 -588
rect -791 588 -757 604
rect -791 -604 -757 -588
rect -533 588 -499 604
rect -533 -604 -499 -588
rect -275 588 -241 604
rect -275 -604 -241 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 241 588 275 604
rect 241 -604 275 -588
rect 499 588 533 604
rect 499 -604 533 -588
rect 757 588 791 604
rect 757 -604 791 -588
rect 1015 588 1049 604
rect 1015 -604 1049 -588
rect 1273 588 1307 604
rect 1273 -604 1307 -588
rect -1261 -681 -1245 -647
rect -1077 -681 -1061 -647
rect -1003 -681 -987 -647
rect -819 -681 -803 -647
rect -745 -681 -729 -647
rect -561 -681 -545 -647
rect -487 -681 -471 -647
rect -303 -681 -287 -647
rect -229 -681 -213 -647
rect -45 -681 -29 -647
rect 29 -681 45 -647
rect 213 -681 229 -647
rect 287 -681 303 -647
rect 471 -681 487 -647
rect 545 -681 561 -647
rect 729 -681 745 -647
rect 803 -681 819 -647
rect 987 -681 1003 -647
rect 1061 -681 1077 -647
rect 1245 -681 1261 -647
rect -1421 -749 -1387 -687
rect 1387 -749 1421 -687
rect -1421 -783 -1325 -749
rect 1325 -783 1421 -749
<< viali >>
rect -1245 647 -1077 681
rect -987 647 -819 681
rect -729 647 -561 681
rect -471 647 -303 681
rect -213 647 -45 681
rect 45 647 213 681
rect 303 647 471 681
rect 561 647 729 681
rect 819 647 987 681
rect 1077 647 1245 681
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect -1245 -681 -1077 -647
rect -987 -681 -819 -647
rect -729 -681 -561 -647
rect -471 -681 -303 -647
rect -213 -681 -45 -647
rect 45 -681 213 -647
rect 303 -681 471 -647
rect 561 -681 729 -647
rect 819 -681 987 -647
rect 1077 -681 1245 -647
<< metal1 >>
rect -1257 681 -1065 687
rect -1257 647 -1245 681
rect -1077 647 -1065 681
rect -1257 641 -1065 647
rect -999 681 -807 687
rect -999 647 -987 681
rect -819 647 -807 681
rect -999 641 -807 647
rect -741 681 -549 687
rect -741 647 -729 681
rect -561 647 -549 681
rect -741 641 -549 647
rect -483 681 -291 687
rect -483 647 -471 681
rect -303 647 -291 681
rect -483 641 -291 647
rect -225 681 -33 687
rect -225 647 -213 681
rect -45 647 -33 681
rect -225 641 -33 647
rect 33 681 225 687
rect 33 647 45 681
rect 213 647 225 681
rect 33 641 225 647
rect 291 681 483 687
rect 291 647 303 681
rect 471 647 483 681
rect 291 641 483 647
rect 549 681 741 687
rect 549 647 561 681
rect 729 647 741 681
rect 549 641 741 647
rect 807 681 999 687
rect 807 647 819 681
rect 987 647 999 681
rect 807 641 999 647
rect 1065 681 1257 687
rect 1065 647 1077 681
rect 1245 647 1257 681
rect 1065 641 1257 647
rect -1313 588 -1267 600
rect -1313 -588 -1307 588
rect -1273 -588 -1267 588
rect -1313 -600 -1267 -588
rect -1055 588 -1009 600
rect -1055 -588 -1049 588
rect -1015 -588 -1009 588
rect -1055 -600 -1009 -588
rect -797 588 -751 600
rect -797 -588 -791 588
rect -757 -588 -751 588
rect -797 -600 -751 -588
rect -539 588 -493 600
rect -539 -588 -533 588
rect -499 -588 -493 588
rect -539 -600 -493 -588
rect -281 588 -235 600
rect -281 -588 -275 588
rect -241 -588 -235 588
rect -281 -600 -235 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 235 588 281 600
rect 235 -588 241 588
rect 275 -588 281 588
rect 235 -600 281 -588
rect 493 588 539 600
rect 493 -588 499 588
rect 533 -588 539 588
rect 493 -600 539 -588
rect 751 588 797 600
rect 751 -588 757 588
rect 791 -588 797 588
rect 751 -600 797 -588
rect 1009 588 1055 600
rect 1009 -588 1015 588
rect 1049 -588 1055 588
rect 1009 -600 1055 -588
rect 1267 588 1313 600
rect 1267 -588 1273 588
rect 1307 -588 1313 588
rect 1267 -600 1313 -588
rect -1257 -647 -1065 -641
rect -1257 -681 -1245 -647
rect -1077 -681 -1065 -647
rect -1257 -687 -1065 -681
rect -999 -647 -807 -641
rect -999 -681 -987 -647
rect -819 -681 -807 -647
rect -999 -687 -807 -681
rect -741 -647 -549 -641
rect -741 -681 -729 -647
rect -561 -681 -549 -647
rect -741 -687 -549 -681
rect -483 -647 -291 -641
rect -483 -681 -471 -647
rect -303 -681 -291 -647
rect -483 -687 -291 -681
rect -225 -647 -33 -641
rect -225 -681 -213 -647
rect -45 -681 -33 -647
rect -225 -687 -33 -681
rect 33 -647 225 -641
rect 33 -681 45 -647
rect 213 -681 225 -647
rect 33 -687 225 -681
rect 291 -647 483 -641
rect 291 -681 303 -647
rect 471 -681 483 -647
rect 291 -687 483 -681
rect 549 -647 741 -641
rect 549 -681 561 -647
rect 729 -681 741 -647
rect 549 -687 741 -681
rect 807 -647 999 -641
rect 807 -681 819 -647
rect 987 -681 999 -647
rect 807 -687 999 -681
rect 1065 -647 1257 -641
rect 1065 -681 1077 -647
rect 1245 -681 1257 -647
rect 1065 -687 1257 -681
<< properties >>
string FIXED_BBOX -1404 -766 1404 766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
