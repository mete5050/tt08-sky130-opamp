magic
tech sky130B
magscale 1 2
timestamp 1768735072
<< error_p >>
rect -3510 681 -3452 687
rect -3392 681 -3334 687
rect -3274 681 -3216 687
rect -3156 681 -3098 687
rect -3038 681 -2980 687
rect -2920 681 -2862 687
rect -2802 681 -2744 687
rect -2684 681 -2626 687
rect -2566 681 -2508 687
rect -2448 681 -2390 687
rect -2330 681 -2272 687
rect -2212 681 -2154 687
rect -2094 681 -2036 687
rect -1976 681 -1918 687
rect -1858 681 -1800 687
rect -1740 681 -1682 687
rect -1622 681 -1564 687
rect -1504 681 -1446 687
rect -1386 681 -1328 687
rect -1268 681 -1210 687
rect -1150 681 -1092 687
rect -1032 681 -974 687
rect -914 681 -856 687
rect -796 681 -738 687
rect -678 681 -620 687
rect -560 681 -502 687
rect -442 681 -384 687
rect -324 681 -266 687
rect -206 681 -148 687
rect -88 681 -30 687
rect 30 681 88 687
rect 148 681 206 687
rect 266 681 324 687
rect 384 681 442 687
rect 502 681 560 687
rect 620 681 678 687
rect 738 681 796 687
rect 856 681 914 687
rect 974 681 1032 687
rect 1092 681 1150 687
rect 1210 681 1268 687
rect 1328 681 1386 687
rect 1446 681 1504 687
rect 1564 681 1622 687
rect 1682 681 1740 687
rect 1800 681 1858 687
rect 1918 681 1976 687
rect 2036 681 2094 687
rect 2154 681 2212 687
rect 2272 681 2330 687
rect 2390 681 2448 687
rect 2508 681 2566 687
rect 2626 681 2684 687
rect 2744 681 2802 687
rect 2862 681 2920 687
rect 2980 681 3038 687
rect 3098 681 3156 687
rect 3216 681 3274 687
rect 3334 681 3392 687
rect 3452 681 3510 687
rect -3510 647 -3498 681
rect -3392 647 -3380 681
rect -3274 647 -3262 681
rect -3156 647 -3144 681
rect -3038 647 -3026 681
rect -2920 647 -2908 681
rect -2802 647 -2790 681
rect -2684 647 -2672 681
rect -2566 647 -2554 681
rect -2448 647 -2436 681
rect -2330 647 -2318 681
rect -2212 647 -2200 681
rect -2094 647 -2082 681
rect -1976 647 -1964 681
rect -1858 647 -1846 681
rect -1740 647 -1728 681
rect -1622 647 -1610 681
rect -1504 647 -1492 681
rect -1386 647 -1374 681
rect -1268 647 -1256 681
rect -1150 647 -1138 681
rect -1032 647 -1020 681
rect -914 647 -902 681
rect -796 647 -784 681
rect -678 647 -666 681
rect -560 647 -548 681
rect -442 647 -430 681
rect -324 647 -312 681
rect -206 647 -194 681
rect -88 647 -76 681
rect 30 647 42 681
rect 148 647 160 681
rect 266 647 278 681
rect 384 647 396 681
rect 502 647 514 681
rect 620 647 632 681
rect 738 647 750 681
rect 856 647 868 681
rect 974 647 986 681
rect 1092 647 1104 681
rect 1210 647 1222 681
rect 1328 647 1340 681
rect 1446 647 1458 681
rect 1564 647 1576 681
rect 1682 647 1694 681
rect 1800 647 1812 681
rect 1918 647 1930 681
rect 2036 647 2048 681
rect 2154 647 2166 681
rect 2272 647 2284 681
rect 2390 647 2402 681
rect 2508 647 2520 681
rect 2626 647 2638 681
rect 2744 647 2756 681
rect 2862 647 2874 681
rect 2980 647 2992 681
rect 3098 647 3110 681
rect 3216 647 3228 681
rect 3334 647 3346 681
rect 3452 647 3464 681
rect -3510 641 -3452 647
rect -3392 641 -3334 647
rect -3274 641 -3216 647
rect -3156 641 -3098 647
rect -3038 641 -2980 647
rect -2920 641 -2862 647
rect -2802 641 -2744 647
rect -2684 641 -2626 647
rect -2566 641 -2508 647
rect -2448 641 -2390 647
rect -2330 641 -2272 647
rect -2212 641 -2154 647
rect -2094 641 -2036 647
rect -1976 641 -1918 647
rect -1858 641 -1800 647
rect -1740 641 -1682 647
rect -1622 641 -1564 647
rect -1504 641 -1446 647
rect -1386 641 -1328 647
rect -1268 641 -1210 647
rect -1150 641 -1092 647
rect -1032 641 -974 647
rect -914 641 -856 647
rect -796 641 -738 647
rect -678 641 -620 647
rect -560 641 -502 647
rect -442 641 -384 647
rect -324 641 -266 647
rect -206 641 -148 647
rect -88 641 -30 647
rect 30 641 88 647
rect 148 641 206 647
rect 266 641 324 647
rect 384 641 442 647
rect 502 641 560 647
rect 620 641 678 647
rect 738 641 796 647
rect 856 641 914 647
rect 974 641 1032 647
rect 1092 641 1150 647
rect 1210 641 1268 647
rect 1328 641 1386 647
rect 1446 641 1504 647
rect 1564 641 1622 647
rect 1682 641 1740 647
rect 1800 641 1858 647
rect 1918 641 1976 647
rect 2036 641 2094 647
rect 2154 641 2212 647
rect 2272 641 2330 647
rect 2390 641 2448 647
rect 2508 641 2566 647
rect 2626 641 2684 647
rect 2744 641 2802 647
rect 2862 641 2920 647
rect 2980 641 3038 647
rect 3098 641 3156 647
rect 3216 641 3274 647
rect 3334 641 3392 647
rect 3452 641 3510 647
rect -3510 -647 -3452 -641
rect -3392 -647 -3334 -641
rect -3274 -647 -3216 -641
rect -3156 -647 -3098 -641
rect -3038 -647 -2980 -641
rect -2920 -647 -2862 -641
rect -2802 -647 -2744 -641
rect -2684 -647 -2626 -641
rect -2566 -647 -2508 -641
rect -2448 -647 -2390 -641
rect -2330 -647 -2272 -641
rect -2212 -647 -2154 -641
rect -2094 -647 -2036 -641
rect -1976 -647 -1918 -641
rect -1858 -647 -1800 -641
rect -1740 -647 -1682 -641
rect -1622 -647 -1564 -641
rect -1504 -647 -1446 -641
rect -1386 -647 -1328 -641
rect -1268 -647 -1210 -641
rect -1150 -647 -1092 -641
rect -1032 -647 -974 -641
rect -914 -647 -856 -641
rect -796 -647 -738 -641
rect -678 -647 -620 -641
rect -560 -647 -502 -641
rect -442 -647 -384 -641
rect -324 -647 -266 -641
rect -206 -647 -148 -641
rect -88 -647 -30 -641
rect 30 -647 88 -641
rect 148 -647 206 -641
rect 266 -647 324 -641
rect 384 -647 442 -641
rect 502 -647 560 -641
rect 620 -647 678 -641
rect 738 -647 796 -641
rect 856 -647 914 -641
rect 974 -647 1032 -641
rect 1092 -647 1150 -641
rect 1210 -647 1268 -641
rect 1328 -647 1386 -641
rect 1446 -647 1504 -641
rect 1564 -647 1622 -641
rect 1682 -647 1740 -641
rect 1800 -647 1858 -641
rect 1918 -647 1976 -641
rect 2036 -647 2094 -641
rect 2154 -647 2212 -641
rect 2272 -647 2330 -641
rect 2390 -647 2448 -641
rect 2508 -647 2566 -641
rect 2626 -647 2684 -641
rect 2744 -647 2802 -641
rect 2862 -647 2920 -641
rect 2980 -647 3038 -641
rect 3098 -647 3156 -641
rect 3216 -647 3274 -641
rect 3334 -647 3392 -641
rect 3452 -647 3510 -641
rect -3510 -681 -3498 -647
rect -3392 -681 -3380 -647
rect -3274 -681 -3262 -647
rect -3156 -681 -3144 -647
rect -3038 -681 -3026 -647
rect -2920 -681 -2908 -647
rect -2802 -681 -2790 -647
rect -2684 -681 -2672 -647
rect -2566 -681 -2554 -647
rect -2448 -681 -2436 -647
rect -2330 -681 -2318 -647
rect -2212 -681 -2200 -647
rect -2094 -681 -2082 -647
rect -1976 -681 -1964 -647
rect -1858 -681 -1846 -647
rect -1740 -681 -1728 -647
rect -1622 -681 -1610 -647
rect -1504 -681 -1492 -647
rect -1386 -681 -1374 -647
rect -1268 -681 -1256 -647
rect -1150 -681 -1138 -647
rect -1032 -681 -1020 -647
rect -914 -681 -902 -647
rect -796 -681 -784 -647
rect -678 -681 -666 -647
rect -560 -681 -548 -647
rect -442 -681 -430 -647
rect -324 -681 -312 -647
rect -206 -681 -194 -647
rect -88 -681 -76 -647
rect 30 -681 42 -647
rect 148 -681 160 -647
rect 266 -681 278 -647
rect 384 -681 396 -647
rect 502 -681 514 -647
rect 620 -681 632 -647
rect 738 -681 750 -647
rect 856 -681 868 -647
rect 974 -681 986 -647
rect 1092 -681 1104 -647
rect 1210 -681 1222 -647
rect 1328 -681 1340 -647
rect 1446 -681 1458 -647
rect 1564 -681 1576 -647
rect 1682 -681 1694 -647
rect 1800 -681 1812 -647
rect 1918 -681 1930 -647
rect 2036 -681 2048 -647
rect 2154 -681 2166 -647
rect 2272 -681 2284 -647
rect 2390 -681 2402 -647
rect 2508 -681 2520 -647
rect 2626 -681 2638 -647
rect 2744 -681 2756 -647
rect 2862 -681 2874 -647
rect 2980 -681 2992 -647
rect 3098 -681 3110 -647
rect 3216 -681 3228 -647
rect 3334 -681 3346 -647
rect 3452 -681 3464 -647
rect -3510 -687 -3452 -681
rect -3392 -687 -3334 -681
rect -3274 -687 -3216 -681
rect -3156 -687 -3098 -681
rect -3038 -687 -2980 -681
rect -2920 -687 -2862 -681
rect -2802 -687 -2744 -681
rect -2684 -687 -2626 -681
rect -2566 -687 -2508 -681
rect -2448 -687 -2390 -681
rect -2330 -687 -2272 -681
rect -2212 -687 -2154 -681
rect -2094 -687 -2036 -681
rect -1976 -687 -1918 -681
rect -1858 -687 -1800 -681
rect -1740 -687 -1682 -681
rect -1622 -687 -1564 -681
rect -1504 -687 -1446 -681
rect -1386 -687 -1328 -681
rect -1268 -687 -1210 -681
rect -1150 -687 -1092 -681
rect -1032 -687 -974 -681
rect -914 -687 -856 -681
rect -796 -687 -738 -681
rect -678 -687 -620 -681
rect -560 -687 -502 -681
rect -442 -687 -384 -681
rect -324 -687 -266 -681
rect -206 -687 -148 -681
rect -88 -687 -30 -681
rect 30 -687 88 -681
rect 148 -687 206 -681
rect 266 -687 324 -681
rect 384 -687 442 -681
rect 502 -687 560 -681
rect 620 -687 678 -681
rect 738 -687 796 -681
rect 856 -687 914 -681
rect 974 -687 1032 -681
rect 1092 -687 1150 -681
rect 1210 -687 1268 -681
rect 1328 -687 1386 -681
rect 1446 -687 1504 -681
rect 1564 -687 1622 -681
rect 1682 -687 1740 -681
rect 1800 -687 1858 -681
rect 1918 -687 1976 -681
rect 2036 -687 2094 -681
rect 2154 -687 2212 -681
rect 2272 -687 2330 -681
rect 2390 -687 2448 -681
rect 2508 -687 2566 -681
rect 2626 -687 2684 -681
rect 2744 -687 2802 -681
rect 2862 -687 2920 -681
rect 2980 -687 3038 -681
rect 3098 -687 3156 -681
rect 3216 -687 3274 -681
rect 3334 -687 3392 -681
rect 3452 -687 3510 -681
<< nwell >>
rect -3605 -700 3605 700
<< pmos >>
rect -3511 -600 -3451 600
rect -3393 -600 -3333 600
rect -3275 -600 -3215 600
rect -3157 -600 -3097 600
rect -3039 -600 -2979 600
rect -2921 -600 -2861 600
rect -2803 -600 -2743 600
rect -2685 -600 -2625 600
rect -2567 -600 -2507 600
rect -2449 -600 -2389 600
rect -2331 -600 -2271 600
rect -2213 -600 -2153 600
rect -2095 -600 -2035 600
rect -1977 -600 -1917 600
rect -1859 -600 -1799 600
rect -1741 -600 -1681 600
rect -1623 -600 -1563 600
rect -1505 -600 -1445 600
rect -1387 -600 -1327 600
rect -1269 -600 -1209 600
rect -1151 -600 -1091 600
rect -1033 -600 -973 600
rect -915 -600 -855 600
rect -797 -600 -737 600
rect -679 -600 -619 600
rect -561 -600 -501 600
rect -443 -600 -383 600
rect -325 -600 -265 600
rect -207 -600 -147 600
rect -89 -600 -29 600
rect 29 -600 89 600
rect 147 -600 207 600
rect 265 -600 325 600
rect 383 -600 443 600
rect 501 -600 561 600
rect 619 -600 679 600
rect 737 -600 797 600
rect 855 -600 915 600
rect 973 -600 1033 600
rect 1091 -600 1151 600
rect 1209 -600 1269 600
rect 1327 -600 1387 600
rect 1445 -600 1505 600
rect 1563 -600 1623 600
rect 1681 -600 1741 600
rect 1799 -600 1859 600
rect 1917 -600 1977 600
rect 2035 -600 2095 600
rect 2153 -600 2213 600
rect 2271 -600 2331 600
rect 2389 -600 2449 600
rect 2507 -600 2567 600
rect 2625 -600 2685 600
rect 2743 -600 2803 600
rect 2861 -600 2921 600
rect 2979 -600 3039 600
rect 3097 -600 3157 600
rect 3215 -600 3275 600
rect 3333 -600 3393 600
rect 3451 -600 3511 600
<< pdiff >>
rect -3569 588 -3511 600
rect -3569 -588 -3557 588
rect -3523 -588 -3511 588
rect -3569 -600 -3511 -588
rect -3451 588 -3393 600
rect -3451 -588 -3439 588
rect -3405 -588 -3393 588
rect -3451 -600 -3393 -588
rect -3333 588 -3275 600
rect -3333 -588 -3321 588
rect -3287 -588 -3275 588
rect -3333 -600 -3275 -588
rect -3215 588 -3157 600
rect -3215 -588 -3203 588
rect -3169 -588 -3157 588
rect -3215 -600 -3157 -588
rect -3097 588 -3039 600
rect -3097 -588 -3085 588
rect -3051 -588 -3039 588
rect -3097 -600 -3039 -588
rect -2979 588 -2921 600
rect -2979 -588 -2967 588
rect -2933 -588 -2921 588
rect -2979 -600 -2921 -588
rect -2861 588 -2803 600
rect -2861 -588 -2849 588
rect -2815 -588 -2803 588
rect -2861 -600 -2803 -588
rect -2743 588 -2685 600
rect -2743 -588 -2731 588
rect -2697 -588 -2685 588
rect -2743 -600 -2685 -588
rect -2625 588 -2567 600
rect -2625 -588 -2613 588
rect -2579 -588 -2567 588
rect -2625 -600 -2567 -588
rect -2507 588 -2449 600
rect -2507 -588 -2495 588
rect -2461 -588 -2449 588
rect -2507 -600 -2449 -588
rect -2389 588 -2331 600
rect -2389 -588 -2377 588
rect -2343 -588 -2331 588
rect -2389 -600 -2331 -588
rect -2271 588 -2213 600
rect -2271 -588 -2259 588
rect -2225 -588 -2213 588
rect -2271 -600 -2213 -588
rect -2153 588 -2095 600
rect -2153 -588 -2141 588
rect -2107 -588 -2095 588
rect -2153 -600 -2095 -588
rect -2035 588 -1977 600
rect -2035 -588 -2023 588
rect -1989 -588 -1977 588
rect -2035 -600 -1977 -588
rect -1917 588 -1859 600
rect -1917 -588 -1905 588
rect -1871 -588 -1859 588
rect -1917 -600 -1859 -588
rect -1799 588 -1741 600
rect -1799 -588 -1787 588
rect -1753 -588 -1741 588
rect -1799 -600 -1741 -588
rect -1681 588 -1623 600
rect -1681 -588 -1669 588
rect -1635 -588 -1623 588
rect -1681 -600 -1623 -588
rect -1563 588 -1505 600
rect -1563 -588 -1551 588
rect -1517 -588 -1505 588
rect -1563 -600 -1505 -588
rect -1445 588 -1387 600
rect -1445 -588 -1433 588
rect -1399 -588 -1387 588
rect -1445 -600 -1387 -588
rect -1327 588 -1269 600
rect -1327 -588 -1315 588
rect -1281 -588 -1269 588
rect -1327 -600 -1269 -588
rect -1209 588 -1151 600
rect -1209 -588 -1197 588
rect -1163 -588 -1151 588
rect -1209 -600 -1151 -588
rect -1091 588 -1033 600
rect -1091 -588 -1079 588
rect -1045 -588 -1033 588
rect -1091 -600 -1033 -588
rect -973 588 -915 600
rect -973 -588 -961 588
rect -927 -588 -915 588
rect -973 -600 -915 -588
rect -855 588 -797 600
rect -855 -588 -843 588
rect -809 -588 -797 588
rect -855 -600 -797 -588
rect -737 588 -679 600
rect -737 -588 -725 588
rect -691 -588 -679 588
rect -737 -600 -679 -588
rect -619 588 -561 600
rect -619 -588 -607 588
rect -573 -588 -561 588
rect -619 -600 -561 -588
rect -501 588 -443 600
rect -501 -588 -489 588
rect -455 -588 -443 588
rect -501 -600 -443 -588
rect -383 588 -325 600
rect -383 -588 -371 588
rect -337 -588 -325 588
rect -383 -600 -325 -588
rect -265 588 -207 600
rect -265 -588 -253 588
rect -219 -588 -207 588
rect -265 -600 -207 -588
rect -147 588 -89 600
rect -147 -588 -135 588
rect -101 -588 -89 588
rect -147 -600 -89 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 89 588 147 600
rect 89 -588 101 588
rect 135 -588 147 588
rect 89 -600 147 -588
rect 207 588 265 600
rect 207 -588 219 588
rect 253 -588 265 588
rect 207 -600 265 -588
rect 325 588 383 600
rect 325 -588 337 588
rect 371 -588 383 588
rect 325 -600 383 -588
rect 443 588 501 600
rect 443 -588 455 588
rect 489 -588 501 588
rect 443 -600 501 -588
rect 561 588 619 600
rect 561 -588 573 588
rect 607 -588 619 588
rect 561 -600 619 -588
rect 679 588 737 600
rect 679 -588 691 588
rect 725 -588 737 588
rect 679 -600 737 -588
rect 797 588 855 600
rect 797 -588 809 588
rect 843 -588 855 588
rect 797 -600 855 -588
rect 915 588 973 600
rect 915 -588 927 588
rect 961 -588 973 588
rect 915 -600 973 -588
rect 1033 588 1091 600
rect 1033 -588 1045 588
rect 1079 -588 1091 588
rect 1033 -600 1091 -588
rect 1151 588 1209 600
rect 1151 -588 1163 588
rect 1197 -588 1209 588
rect 1151 -600 1209 -588
rect 1269 588 1327 600
rect 1269 -588 1281 588
rect 1315 -588 1327 588
rect 1269 -600 1327 -588
rect 1387 588 1445 600
rect 1387 -588 1399 588
rect 1433 -588 1445 588
rect 1387 -600 1445 -588
rect 1505 588 1563 600
rect 1505 -588 1517 588
rect 1551 -588 1563 588
rect 1505 -600 1563 -588
rect 1623 588 1681 600
rect 1623 -588 1635 588
rect 1669 -588 1681 588
rect 1623 -600 1681 -588
rect 1741 588 1799 600
rect 1741 -588 1753 588
rect 1787 -588 1799 588
rect 1741 -600 1799 -588
rect 1859 588 1917 600
rect 1859 -588 1871 588
rect 1905 -588 1917 588
rect 1859 -600 1917 -588
rect 1977 588 2035 600
rect 1977 -588 1989 588
rect 2023 -588 2035 588
rect 1977 -600 2035 -588
rect 2095 588 2153 600
rect 2095 -588 2107 588
rect 2141 -588 2153 588
rect 2095 -600 2153 -588
rect 2213 588 2271 600
rect 2213 -588 2225 588
rect 2259 -588 2271 588
rect 2213 -600 2271 -588
rect 2331 588 2389 600
rect 2331 -588 2343 588
rect 2377 -588 2389 588
rect 2331 -600 2389 -588
rect 2449 588 2507 600
rect 2449 -588 2461 588
rect 2495 -588 2507 588
rect 2449 -600 2507 -588
rect 2567 588 2625 600
rect 2567 -588 2579 588
rect 2613 -588 2625 588
rect 2567 -600 2625 -588
rect 2685 588 2743 600
rect 2685 -588 2697 588
rect 2731 -588 2743 588
rect 2685 -600 2743 -588
rect 2803 588 2861 600
rect 2803 -588 2815 588
rect 2849 -588 2861 588
rect 2803 -600 2861 -588
rect 2921 588 2979 600
rect 2921 -588 2933 588
rect 2967 -588 2979 588
rect 2921 -600 2979 -588
rect 3039 588 3097 600
rect 3039 -588 3051 588
rect 3085 -588 3097 588
rect 3039 -600 3097 -588
rect 3157 588 3215 600
rect 3157 -588 3169 588
rect 3203 -588 3215 588
rect 3157 -600 3215 -588
rect 3275 588 3333 600
rect 3275 -588 3287 588
rect 3321 -588 3333 588
rect 3275 -600 3333 -588
rect 3393 588 3451 600
rect 3393 -588 3405 588
rect 3439 -588 3451 588
rect 3393 -600 3451 -588
rect 3511 588 3569 600
rect 3511 -588 3523 588
rect 3557 -588 3569 588
rect 3511 -600 3569 -588
<< pdiffc >>
rect -3557 -588 -3523 588
rect -3439 -588 -3405 588
rect -3321 -588 -3287 588
rect -3203 -588 -3169 588
rect -3085 -588 -3051 588
rect -2967 -588 -2933 588
rect -2849 -588 -2815 588
rect -2731 -588 -2697 588
rect -2613 -588 -2579 588
rect -2495 -588 -2461 588
rect -2377 -588 -2343 588
rect -2259 -588 -2225 588
rect -2141 -588 -2107 588
rect -2023 -588 -1989 588
rect -1905 -588 -1871 588
rect -1787 -588 -1753 588
rect -1669 -588 -1635 588
rect -1551 -588 -1517 588
rect -1433 -588 -1399 588
rect -1315 -588 -1281 588
rect -1197 -588 -1163 588
rect -1079 -588 -1045 588
rect -961 -588 -927 588
rect -843 -588 -809 588
rect -725 -588 -691 588
rect -607 -588 -573 588
rect -489 -588 -455 588
rect -371 -588 -337 588
rect -253 -588 -219 588
rect -135 -588 -101 588
rect -17 -588 17 588
rect 101 -588 135 588
rect 219 -588 253 588
rect 337 -588 371 588
rect 455 -588 489 588
rect 573 -588 607 588
rect 691 -588 725 588
rect 809 -588 843 588
rect 927 -588 961 588
rect 1045 -588 1079 588
rect 1163 -588 1197 588
rect 1281 -588 1315 588
rect 1399 -588 1433 588
rect 1517 -588 1551 588
rect 1635 -588 1669 588
rect 1753 -588 1787 588
rect 1871 -588 1905 588
rect 1989 -588 2023 588
rect 2107 -588 2141 588
rect 2225 -588 2259 588
rect 2343 -588 2377 588
rect 2461 -588 2495 588
rect 2579 -588 2613 588
rect 2697 -588 2731 588
rect 2815 -588 2849 588
rect 2933 -588 2967 588
rect 3051 -588 3085 588
rect 3169 -588 3203 588
rect 3287 -588 3321 588
rect 3405 -588 3439 588
rect 3523 -588 3557 588
<< poly >>
rect -3514 681 -3448 697
rect -3514 647 -3498 681
rect -3464 647 -3448 681
rect -3514 631 -3448 647
rect -3396 681 -3330 697
rect -3396 647 -3380 681
rect -3346 647 -3330 681
rect -3396 631 -3330 647
rect -3278 681 -3212 697
rect -3278 647 -3262 681
rect -3228 647 -3212 681
rect -3278 631 -3212 647
rect -3160 681 -3094 697
rect -3160 647 -3144 681
rect -3110 647 -3094 681
rect -3160 631 -3094 647
rect -3042 681 -2976 697
rect -3042 647 -3026 681
rect -2992 647 -2976 681
rect -3042 631 -2976 647
rect -2924 681 -2858 697
rect -2924 647 -2908 681
rect -2874 647 -2858 681
rect -2924 631 -2858 647
rect -2806 681 -2740 697
rect -2806 647 -2790 681
rect -2756 647 -2740 681
rect -2806 631 -2740 647
rect -2688 681 -2622 697
rect -2688 647 -2672 681
rect -2638 647 -2622 681
rect -2688 631 -2622 647
rect -2570 681 -2504 697
rect -2570 647 -2554 681
rect -2520 647 -2504 681
rect -2570 631 -2504 647
rect -2452 681 -2386 697
rect -2452 647 -2436 681
rect -2402 647 -2386 681
rect -2452 631 -2386 647
rect -2334 681 -2268 697
rect -2334 647 -2318 681
rect -2284 647 -2268 681
rect -2334 631 -2268 647
rect -2216 681 -2150 697
rect -2216 647 -2200 681
rect -2166 647 -2150 681
rect -2216 631 -2150 647
rect -2098 681 -2032 697
rect -2098 647 -2082 681
rect -2048 647 -2032 681
rect -2098 631 -2032 647
rect -1980 681 -1914 697
rect -1980 647 -1964 681
rect -1930 647 -1914 681
rect -1980 631 -1914 647
rect -1862 681 -1796 697
rect -1862 647 -1846 681
rect -1812 647 -1796 681
rect -1862 631 -1796 647
rect -1744 681 -1678 697
rect -1744 647 -1728 681
rect -1694 647 -1678 681
rect -1744 631 -1678 647
rect -1626 681 -1560 697
rect -1626 647 -1610 681
rect -1576 647 -1560 681
rect -1626 631 -1560 647
rect -1508 681 -1442 697
rect -1508 647 -1492 681
rect -1458 647 -1442 681
rect -1508 631 -1442 647
rect -1390 681 -1324 697
rect -1390 647 -1374 681
rect -1340 647 -1324 681
rect -1390 631 -1324 647
rect -1272 681 -1206 697
rect -1272 647 -1256 681
rect -1222 647 -1206 681
rect -1272 631 -1206 647
rect -1154 681 -1088 697
rect -1154 647 -1138 681
rect -1104 647 -1088 681
rect -1154 631 -1088 647
rect -1036 681 -970 697
rect -1036 647 -1020 681
rect -986 647 -970 681
rect -1036 631 -970 647
rect -918 681 -852 697
rect -918 647 -902 681
rect -868 647 -852 681
rect -918 631 -852 647
rect -800 681 -734 697
rect -800 647 -784 681
rect -750 647 -734 681
rect -800 631 -734 647
rect -682 681 -616 697
rect -682 647 -666 681
rect -632 647 -616 681
rect -682 631 -616 647
rect -564 681 -498 697
rect -564 647 -548 681
rect -514 647 -498 681
rect -564 631 -498 647
rect -446 681 -380 697
rect -446 647 -430 681
rect -396 647 -380 681
rect -446 631 -380 647
rect -328 681 -262 697
rect -328 647 -312 681
rect -278 647 -262 681
rect -328 631 -262 647
rect -210 681 -144 697
rect -210 647 -194 681
rect -160 647 -144 681
rect -210 631 -144 647
rect -92 681 -26 697
rect -92 647 -76 681
rect -42 647 -26 681
rect -92 631 -26 647
rect 26 681 92 697
rect 26 647 42 681
rect 76 647 92 681
rect 26 631 92 647
rect 144 681 210 697
rect 144 647 160 681
rect 194 647 210 681
rect 144 631 210 647
rect 262 681 328 697
rect 262 647 278 681
rect 312 647 328 681
rect 262 631 328 647
rect 380 681 446 697
rect 380 647 396 681
rect 430 647 446 681
rect 380 631 446 647
rect 498 681 564 697
rect 498 647 514 681
rect 548 647 564 681
rect 498 631 564 647
rect 616 681 682 697
rect 616 647 632 681
rect 666 647 682 681
rect 616 631 682 647
rect 734 681 800 697
rect 734 647 750 681
rect 784 647 800 681
rect 734 631 800 647
rect 852 681 918 697
rect 852 647 868 681
rect 902 647 918 681
rect 852 631 918 647
rect 970 681 1036 697
rect 970 647 986 681
rect 1020 647 1036 681
rect 970 631 1036 647
rect 1088 681 1154 697
rect 1088 647 1104 681
rect 1138 647 1154 681
rect 1088 631 1154 647
rect 1206 681 1272 697
rect 1206 647 1222 681
rect 1256 647 1272 681
rect 1206 631 1272 647
rect 1324 681 1390 697
rect 1324 647 1340 681
rect 1374 647 1390 681
rect 1324 631 1390 647
rect 1442 681 1508 697
rect 1442 647 1458 681
rect 1492 647 1508 681
rect 1442 631 1508 647
rect 1560 681 1626 697
rect 1560 647 1576 681
rect 1610 647 1626 681
rect 1560 631 1626 647
rect 1678 681 1744 697
rect 1678 647 1694 681
rect 1728 647 1744 681
rect 1678 631 1744 647
rect 1796 681 1862 697
rect 1796 647 1812 681
rect 1846 647 1862 681
rect 1796 631 1862 647
rect 1914 681 1980 697
rect 1914 647 1930 681
rect 1964 647 1980 681
rect 1914 631 1980 647
rect 2032 681 2098 697
rect 2032 647 2048 681
rect 2082 647 2098 681
rect 2032 631 2098 647
rect 2150 681 2216 697
rect 2150 647 2166 681
rect 2200 647 2216 681
rect 2150 631 2216 647
rect 2268 681 2334 697
rect 2268 647 2284 681
rect 2318 647 2334 681
rect 2268 631 2334 647
rect 2386 681 2452 697
rect 2386 647 2402 681
rect 2436 647 2452 681
rect 2386 631 2452 647
rect 2504 681 2570 697
rect 2504 647 2520 681
rect 2554 647 2570 681
rect 2504 631 2570 647
rect 2622 681 2688 697
rect 2622 647 2638 681
rect 2672 647 2688 681
rect 2622 631 2688 647
rect 2740 681 2806 697
rect 2740 647 2756 681
rect 2790 647 2806 681
rect 2740 631 2806 647
rect 2858 681 2924 697
rect 2858 647 2874 681
rect 2908 647 2924 681
rect 2858 631 2924 647
rect 2976 681 3042 697
rect 2976 647 2992 681
rect 3026 647 3042 681
rect 2976 631 3042 647
rect 3094 681 3160 697
rect 3094 647 3110 681
rect 3144 647 3160 681
rect 3094 631 3160 647
rect 3212 681 3278 697
rect 3212 647 3228 681
rect 3262 647 3278 681
rect 3212 631 3278 647
rect 3330 681 3396 697
rect 3330 647 3346 681
rect 3380 647 3396 681
rect 3330 631 3396 647
rect 3448 681 3514 697
rect 3448 647 3464 681
rect 3498 647 3514 681
rect 3448 631 3514 647
rect -3511 600 -3451 631
rect -3393 600 -3333 631
rect -3275 600 -3215 631
rect -3157 600 -3097 631
rect -3039 600 -2979 631
rect -2921 600 -2861 631
rect -2803 600 -2743 631
rect -2685 600 -2625 631
rect -2567 600 -2507 631
rect -2449 600 -2389 631
rect -2331 600 -2271 631
rect -2213 600 -2153 631
rect -2095 600 -2035 631
rect -1977 600 -1917 631
rect -1859 600 -1799 631
rect -1741 600 -1681 631
rect -1623 600 -1563 631
rect -1505 600 -1445 631
rect -1387 600 -1327 631
rect -1269 600 -1209 631
rect -1151 600 -1091 631
rect -1033 600 -973 631
rect -915 600 -855 631
rect -797 600 -737 631
rect -679 600 -619 631
rect -561 600 -501 631
rect -443 600 -383 631
rect -325 600 -265 631
rect -207 600 -147 631
rect -89 600 -29 631
rect 29 600 89 631
rect 147 600 207 631
rect 265 600 325 631
rect 383 600 443 631
rect 501 600 561 631
rect 619 600 679 631
rect 737 600 797 631
rect 855 600 915 631
rect 973 600 1033 631
rect 1091 600 1151 631
rect 1209 600 1269 631
rect 1327 600 1387 631
rect 1445 600 1505 631
rect 1563 600 1623 631
rect 1681 600 1741 631
rect 1799 600 1859 631
rect 1917 600 1977 631
rect 2035 600 2095 631
rect 2153 600 2213 631
rect 2271 600 2331 631
rect 2389 600 2449 631
rect 2507 600 2567 631
rect 2625 600 2685 631
rect 2743 600 2803 631
rect 2861 600 2921 631
rect 2979 600 3039 631
rect 3097 600 3157 631
rect 3215 600 3275 631
rect 3333 600 3393 631
rect 3451 600 3511 631
rect -3511 -631 -3451 -600
rect -3393 -631 -3333 -600
rect -3275 -631 -3215 -600
rect -3157 -631 -3097 -600
rect -3039 -631 -2979 -600
rect -2921 -631 -2861 -600
rect -2803 -631 -2743 -600
rect -2685 -631 -2625 -600
rect -2567 -631 -2507 -600
rect -2449 -631 -2389 -600
rect -2331 -631 -2271 -600
rect -2213 -631 -2153 -600
rect -2095 -631 -2035 -600
rect -1977 -631 -1917 -600
rect -1859 -631 -1799 -600
rect -1741 -631 -1681 -600
rect -1623 -631 -1563 -600
rect -1505 -631 -1445 -600
rect -1387 -631 -1327 -600
rect -1269 -631 -1209 -600
rect -1151 -631 -1091 -600
rect -1033 -631 -973 -600
rect -915 -631 -855 -600
rect -797 -631 -737 -600
rect -679 -631 -619 -600
rect -561 -631 -501 -600
rect -443 -631 -383 -600
rect -325 -631 -265 -600
rect -207 -631 -147 -600
rect -89 -631 -29 -600
rect 29 -631 89 -600
rect 147 -631 207 -600
rect 265 -631 325 -600
rect 383 -631 443 -600
rect 501 -631 561 -600
rect 619 -631 679 -600
rect 737 -631 797 -600
rect 855 -631 915 -600
rect 973 -631 1033 -600
rect 1091 -631 1151 -600
rect 1209 -631 1269 -600
rect 1327 -631 1387 -600
rect 1445 -631 1505 -600
rect 1563 -631 1623 -600
rect 1681 -631 1741 -600
rect 1799 -631 1859 -600
rect 1917 -631 1977 -600
rect 2035 -631 2095 -600
rect 2153 -631 2213 -600
rect 2271 -631 2331 -600
rect 2389 -631 2449 -600
rect 2507 -631 2567 -600
rect 2625 -631 2685 -600
rect 2743 -631 2803 -600
rect 2861 -631 2921 -600
rect 2979 -631 3039 -600
rect 3097 -631 3157 -600
rect 3215 -631 3275 -600
rect 3333 -631 3393 -600
rect 3451 -631 3511 -600
rect -3514 -647 -3448 -631
rect -3514 -681 -3498 -647
rect -3464 -681 -3448 -647
rect -3514 -697 -3448 -681
rect -3396 -647 -3330 -631
rect -3396 -681 -3380 -647
rect -3346 -681 -3330 -647
rect -3396 -697 -3330 -681
rect -3278 -647 -3212 -631
rect -3278 -681 -3262 -647
rect -3228 -681 -3212 -647
rect -3278 -697 -3212 -681
rect -3160 -647 -3094 -631
rect -3160 -681 -3144 -647
rect -3110 -681 -3094 -647
rect -3160 -697 -3094 -681
rect -3042 -647 -2976 -631
rect -3042 -681 -3026 -647
rect -2992 -681 -2976 -647
rect -3042 -697 -2976 -681
rect -2924 -647 -2858 -631
rect -2924 -681 -2908 -647
rect -2874 -681 -2858 -647
rect -2924 -697 -2858 -681
rect -2806 -647 -2740 -631
rect -2806 -681 -2790 -647
rect -2756 -681 -2740 -647
rect -2806 -697 -2740 -681
rect -2688 -647 -2622 -631
rect -2688 -681 -2672 -647
rect -2638 -681 -2622 -647
rect -2688 -697 -2622 -681
rect -2570 -647 -2504 -631
rect -2570 -681 -2554 -647
rect -2520 -681 -2504 -647
rect -2570 -697 -2504 -681
rect -2452 -647 -2386 -631
rect -2452 -681 -2436 -647
rect -2402 -681 -2386 -647
rect -2452 -697 -2386 -681
rect -2334 -647 -2268 -631
rect -2334 -681 -2318 -647
rect -2284 -681 -2268 -647
rect -2334 -697 -2268 -681
rect -2216 -647 -2150 -631
rect -2216 -681 -2200 -647
rect -2166 -681 -2150 -647
rect -2216 -697 -2150 -681
rect -2098 -647 -2032 -631
rect -2098 -681 -2082 -647
rect -2048 -681 -2032 -647
rect -2098 -697 -2032 -681
rect -1980 -647 -1914 -631
rect -1980 -681 -1964 -647
rect -1930 -681 -1914 -647
rect -1980 -697 -1914 -681
rect -1862 -647 -1796 -631
rect -1862 -681 -1846 -647
rect -1812 -681 -1796 -647
rect -1862 -697 -1796 -681
rect -1744 -647 -1678 -631
rect -1744 -681 -1728 -647
rect -1694 -681 -1678 -647
rect -1744 -697 -1678 -681
rect -1626 -647 -1560 -631
rect -1626 -681 -1610 -647
rect -1576 -681 -1560 -647
rect -1626 -697 -1560 -681
rect -1508 -647 -1442 -631
rect -1508 -681 -1492 -647
rect -1458 -681 -1442 -647
rect -1508 -697 -1442 -681
rect -1390 -647 -1324 -631
rect -1390 -681 -1374 -647
rect -1340 -681 -1324 -647
rect -1390 -697 -1324 -681
rect -1272 -647 -1206 -631
rect -1272 -681 -1256 -647
rect -1222 -681 -1206 -647
rect -1272 -697 -1206 -681
rect -1154 -647 -1088 -631
rect -1154 -681 -1138 -647
rect -1104 -681 -1088 -647
rect -1154 -697 -1088 -681
rect -1036 -647 -970 -631
rect -1036 -681 -1020 -647
rect -986 -681 -970 -647
rect -1036 -697 -970 -681
rect -918 -647 -852 -631
rect -918 -681 -902 -647
rect -868 -681 -852 -647
rect -918 -697 -852 -681
rect -800 -647 -734 -631
rect -800 -681 -784 -647
rect -750 -681 -734 -647
rect -800 -697 -734 -681
rect -682 -647 -616 -631
rect -682 -681 -666 -647
rect -632 -681 -616 -647
rect -682 -697 -616 -681
rect -564 -647 -498 -631
rect -564 -681 -548 -647
rect -514 -681 -498 -647
rect -564 -697 -498 -681
rect -446 -647 -380 -631
rect -446 -681 -430 -647
rect -396 -681 -380 -647
rect -446 -697 -380 -681
rect -328 -647 -262 -631
rect -328 -681 -312 -647
rect -278 -681 -262 -647
rect -328 -697 -262 -681
rect -210 -647 -144 -631
rect -210 -681 -194 -647
rect -160 -681 -144 -647
rect -210 -697 -144 -681
rect -92 -647 -26 -631
rect -92 -681 -76 -647
rect -42 -681 -26 -647
rect -92 -697 -26 -681
rect 26 -647 92 -631
rect 26 -681 42 -647
rect 76 -681 92 -647
rect 26 -697 92 -681
rect 144 -647 210 -631
rect 144 -681 160 -647
rect 194 -681 210 -647
rect 144 -697 210 -681
rect 262 -647 328 -631
rect 262 -681 278 -647
rect 312 -681 328 -647
rect 262 -697 328 -681
rect 380 -647 446 -631
rect 380 -681 396 -647
rect 430 -681 446 -647
rect 380 -697 446 -681
rect 498 -647 564 -631
rect 498 -681 514 -647
rect 548 -681 564 -647
rect 498 -697 564 -681
rect 616 -647 682 -631
rect 616 -681 632 -647
rect 666 -681 682 -647
rect 616 -697 682 -681
rect 734 -647 800 -631
rect 734 -681 750 -647
rect 784 -681 800 -647
rect 734 -697 800 -681
rect 852 -647 918 -631
rect 852 -681 868 -647
rect 902 -681 918 -647
rect 852 -697 918 -681
rect 970 -647 1036 -631
rect 970 -681 986 -647
rect 1020 -681 1036 -647
rect 970 -697 1036 -681
rect 1088 -647 1154 -631
rect 1088 -681 1104 -647
rect 1138 -681 1154 -647
rect 1088 -697 1154 -681
rect 1206 -647 1272 -631
rect 1206 -681 1222 -647
rect 1256 -681 1272 -647
rect 1206 -697 1272 -681
rect 1324 -647 1390 -631
rect 1324 -681 1340 -647
rect 1374 -681 1390 -647
rect 1324 -697 1390 -681
rect 1442 -647 1508 -631
rect 1442 -681 1458 -647
rect 1492 -681 1508 -647
rect 1442 -697 1508 -681
rect 1560 -647 1626 -631
rect 1560 -681 1576 -647
rect 1610 -681 1626 -647
rect 1560 -697 1626 -681
rect 1678 -647 1744 -631
rect 1678 -681 1694 -647
rect 1728 -681 1744 -647
rect 1678 -697 1744 -681
rect 1796 -647 1862 -631
rect 1796 -681 1812 -647
rect 1846 -681 1862 -647
rect 1796 -697 1862 -681
rect 1914 -647 1980 -631
rect 1914 -681 1930 -647
rect 1964 -681 1980 -647
rect 1914 -697 1980 -681
rect 2032 -647 2098 -631
rect 2032 -681 2048 -647
rect 2082 -681 2098 -647
rect 2032 -697 2098 -681
rect 2150 -647 2216 -631
rect 2150 -681 2166 -647
rect 2200 -681 2216 -647
rect 2150 -697 2216 -681
rect 2268 -647 2334 -631
rect 2268 -681 2284 -647
rect 2318 -681 2334 -647
rect 2268 -697 2334 -681
rect 2386 -647 2452 -631
rect 2386 -681 2402 -647
rect 2436 -681 2452 -647
rect 2386 -697 2452 -681
rect 2504 -647 2570 -631
rect 2504 -681 2520 -647
rect 2554 -681 2570 -647
rect 2504 -697 2570 -681
rect 2622 -647 2688 -631
rect 2622 -681 2638 -647
rect 2672 -681 2688 -647
rect 2622 -697 2688 -681
rect 2740 -647 2806 -631
rect 2740 -681 2756 -647
rect 2790 -681 2806 -647
rect 2740 -697 2806 -681
rect 2858 -647 2924 -631
rect 2858 -681 2874 -647
rect 2908 -681 2924 -647
rect 2858 -697 2924 -681
rect 2976 -647 3042 -631
rect 2976 -681 2992 -647
rect 3026 -681 3042 -647
rect 2976 -697 3042 -681
rect 3094 -647 3160 -631
rect 3094 -681 3110 -647
rect 3144 -681 3160 -647
rect 3094 -697 3160 -681
rect 3212 -647 3278 -631
rect 3212 -681 3228 -647
rect 3262 -681 3278 -647
rect 3212 -697 3278 -681
rect 3330 -647 3396 -631
rect 3330 -681 3346 -647
rect 3380 -681 3396 -647
rect 3330 -697 3396 -681
rect 3448 -647 3514 -631
rect 3448 -681 3464 -647
rect 3498 -681 3514 -647
rect 3448 -697 3514 -681
<< polycont >>
rect -3498 647 -3464 681
rect -3380 647 -3346 681
rect -3262 647 -3228 681
rect -3144 647 -3110 681
rect -3026 647 -2992 681
rect -2908 647 -2874 681
rect -2790 647 -2756 681
rect -2672 647 -2638 681
rect -2554 647 -2520 681
rect -2436 647 -2402 681
rect -2318 647 -2284 681
rect -2200 647 -2166 681
rect -2082 647 -2048 681
rect -1964 647 -1930 681
rect -1846 647 -1812 681
rect -1728 647 -1694 681
rect -1610 647 -1576 681
rect -1492 647 -1458 681
rect -1374 647 -1340 681
rect -1256 647 -1222 681
rect -1138 647 -1104 681
rect -1020 647 -986 681
rect -902 647 -868 681
rect -784 647 -750 681
rect -666 647 -632 681
rect -548 647 -514 681
rect -430 647 -396 681
rect -312 647 -278 681
rect -194 647 -160 681
rect -76 647 -42 681
rect 42 647 76 681
rect 160 647 194 681
rect 278 647 312 681
rect 396 647 430 681
rect 514 647 548 681
rect 632 647 666 681
rect 750 647 784 681
rect 868 647 902 681
rect 986 647 1020 681
rect 1104 647 1138 681
rect 1222 647 1256 681
rect 1340 647 1374 681
rect 1458 647 1492 681
rect 1576 647 1610 681
rect 1694 647 1728 681
rect 1812 647 1846 681
rect 1930 647 1964 681
rect 2048 647 2082 681
rect 2166 647 2200 681
rect 2284 647 2318 681
rect 2402 647 2436 681
rect 2520 647 2554 681
rect 2638 647 2672 681
rect 2756 647 2790 681
rect 2874 647 2908 681
rect 2992 647 3026 681
rect 3110 647 3144 681
rect 3228 647 3262 681
rect 3346 647 3380 681
rect 3464 647 3498 681
rect -3498 -681 -3464 -647
rect -3380 -681 -3346 -647
rect -3262 -681 -3228 -647
rect -3144 -681 -3110 -647
rect -3026 -681 -2992 -647
rect -2908 -681 -2874 -647
rect -2790 -681 -2756 -647
rect -2672 -681 -2638 -647
rect -2554 -681 -2520 -647
rect -2436 -681 -2402 -647
rect -2318 -681 -2284 -647
rect -2200 -681 -2166 -647
rect -2082 -681 -2048 -647
rect -1964 -681 -1930 -647
rect -1846 -681 -1812 -647
rect -1728 -681 -1694 -647
rect -1610 -681 -1576 -647
rect -1492 -681 -1458 -647
rect -1374 -681 -1340 -647
rect -1256 -681 -1222 -647
rect -1138 -681 -1104 -647
rect -1020 -681 -986 -647
rect -902 -681 -868 -647
rect -784 -681 -750 -647
rect -666 -681 -632 -647
rect -548 -681 -514 -647
rect -430 -681 -396 -647
rect -312 -681 -278 -647
rect -194 -681 -160 -647
rect -76 -681 -42 -647
rect 42 -681 76 -647
rect 160 -681 194 -647
rect 278 -681 312 -647
rect 396 -681 430 -647
rect 514 -681 548 -647
rect 632 -681 666 -647
rect 750 -681 784 -647
rect 868 -681 902 -647
rect 986 -681 1020 -647
rect 1104 -681 1138 -647
rect 1222 -681 1256 -647
rect 1340 -681 1374 -647
rect 1458 -681 1492 -647
rect 1576 -681 1610 -647
rect 1694 -681 1728 -647
rect 1812 -681 1846 -647
rect 1930 -681 1964 -647
rect 2048 -681 2082 -647
rect 2166 -681 2200 -647
rect 2284 -681 2318 -647
rect 2402 -681 2436 -647
rect 2520 -681 2554 -647
rect 2638 -681 2672 -647
rect 2756 -681 2790 -647
rect 2874 -681 2908 -647
rect 2992 -681 3026 -647
rect 3110 -681 3144 -647
rect 3228 -681 3262 -647
rect 3346 -681 3380 -647
rect 3464 -681 3498 -647
<< locali >>
rect -3514 647 -3498 681
rect -3464 647 -3448 681
rect -3396 647 -3380 681
rect -3346 647 -3330 681
rect -3278 647 -3262 681
rect -3228 647 -3212 681
rect -3160 647 -3144 681
rect -3110 647 -3094 681
rect -3042 647 -3026 681
rect -2992 647 -2976 681
rect -2924 647 -2908 681
rect -2874 647 -2858 681
rect -2806 647 -2790 681
rect -2756 647 -2740 681
rect -2688 647 -2672 681
rect -2638 647 -2622 681
rect -2570 647 -2554 681
rect -2520 647 -2504 681
rect -2452 647 -2436 681
rect -2402 647 -2386 681
rect -2334 647 -2318 681
rect -2284 647 -2268 681
rect -2216 647 -2200 681
rect -2166 647 -2150 681
rect -2098 647 -2082 681
rect -2048 647 -2032 681
rect -1980 647 -1964 681
rect -1930 647 -1914 681
rect -1862 647 -1846 681
rect -1812 647 -1796 681
rect -1744 647 -1728 681
rect -1694 647 -1678 681
rect -1626 647 -1610 681
rect -1576 647 -1560 681
rect -1508 647 -1492 681
rect -1458 647 -1442 681
rect -1390 647 -1374 681
rect -1340 647 -1324 681
rect -1272 647 -1256 681
rect -1222 647 -1206 681
rect -1154 647 -1138 681
rect -1104 647 -1088 681
rect -1036 647 -1020 681
rect -986 647 -970 681
rect -918 647 -902 681
rect -868 647 -852 681
rect -800 647 -784 681
rect -750 647 -734 681
rect -682 647 -666 681
rect -632 647 -616 681
rect -564 647 -548 681
rect -514 647 -498 681
rect -446 647 -430 681
rect -396 647 -380 681
rect -328 647 -312 681
rect -278 647 -262 681
rect -210 647 -194 681
rect -160 647 -144 681
rect -92 647 -76 681
rect -42 647 -26 681
rect 26 647 42 681
rect 76 647 92 681
rect 144 647 160 681
rect 194 647 210 681
rect 262 647 278 681
rect 312 647 328 681
rect 380 647 396 681
rect 430 647 446 681
rect 498 647 514 681
rect 548 647 564 681
rect 616 647 632 681
rect 666 647 682 681
rect 734 647 750 681
rect 784 647 800 681
rect 852 647 868 681
rect 902 647 918 681
rect 970 647 986 681
rect 1020 647 1036 681
rect 1088 647 1104 681
rect 1138 647 1154 681
rect 1206 647 1222 681
rect 1256 647 1272 681
rect 1324 647 1340 681
rect 1374 647 1390 681
rect 1442 647 1458 681
rect 1492 647 1508 681
rect 1560 647 1576 681
rect 1610 647 1626 681
rect 1678 647 1694 681
rect 1728 647 1744 681
rect 1796 647 1812 681
rect 1846 647 1862 681
rect 1914 647 1930 681
rect 1964 647 1980 681
rect 2032 647 2048 681
rect 2082 647 2098 681
rect 2150 647 2166 681
rect 2200 647 2216 681
rect 2268 647 2284 681
rect 2318 647 2334 681
rect 2386 647 2402 681
rect 2436 647 2452 681
rect 2504 647 2520 681
rect 2554 647 2570 681
rect 2622 647 2638 681
rect 2672 647 2688 681
rect 2740 647 2756 681
rect 2790 647 2806 681
rect 2858 647 2874 681
rect 2908 647 2924 681
rect 2976 647 2992 681
rect 3026 647 3042 681
rect 3094 647 3110 681
rect 3144 647 3160 681
rect 3212 647 3228 681
rect 3262 647 3278 681
rect 3330 647 3346 681
rect 3380 647 3396 681
rect 3448 647 3464 681
rect 3498 647 3514 681
rect -3557 588 -3523 604
rect -3557 -604 -3523 -588
rect -3439 588 -3405 604
rect -3439 -604 -3405 -588
rect -3321 588 -3287 604
rect -3321 -604 -3287 -588
rect -3203 588 -3169 604
rect -3203 -604 -3169 -588
rect -3085 588 -3051 604
rect -3085 -604 -3051 -588
rect -2967 588 -2933 604
rect -2967 -604 -2933 -588
rect -2849 588 -2815 604
rect -2849 -604 -2815 -588
rect -2731 588 -2697 604
rect -2731 -604 -2697 -588
rect -2613 588 -2579 604
rect -2613 -604 -2579 -588
rect -2495 588 -2461 604
rect -2495 -604 -2461 -588
rect -2377 588 -2343 604
rect -2377 -604 -2343 -588
rect -2259 588 -2225 604
rect -2259 -604 -2225 -588
rect -2141 588 -2107 604
rect -2141 -604 -2107 -588
rect -2023 588 -1989 604
rect -2023 -604 -1989 -588
rect -1905 588 -1871 604
rect -1905 -604 -1871 -588
rect -1787 588 -1753 604
rect -1787 -604 -1753 -588
rect -1669 588 -1635 604
rect -1669 -604 -1635 -588
rect -1551 588 -1517 604
rect -1551 -604 -1517 -588
rect -1433 588 -1399 604
rect -1433 -604 -1399 -588
rect -1315 588 -1281 604
rect -1315 -604 -1281 -588
rect -1197 588 -1163 604
rect -1197 -604 -1163 -588
rect -1079 588 -1045 604
rect -1079 -604 -1045 -588
rect -961 588 -927 604
rect -961 -604 -927 -588
rect -843 588 -809 604
rect -843 -604 -809 -588
rect -725 588 -691 604
rect -725 -604 -691 -588
rect -607 588 -573 604
rect -607 -604 -573 -588
rect -489 588 -455 604
rect -489 -604 -455 -588
rect -371 588 -337 604
rect -371 -604 -337 -588
rect -253 588 -219 604
rect -253 -604 -219 -588
rect -135 588 -101 604
rect -135 -604 -101 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 101 588 135 604
rect 101 -604 135 -588
rect 219 588 253 604
rect 219 -604 253 -588
rect 337 588 371 604
rect 337 -604 371 -588
rect 455 588 489 604
rect 455 -604 489 -588
rect 573 588 607 604
rect 573 -604 607 -588
rect 691 588 725 604
rect 691 -604 725 -588
rect 809 588 843 604
rect 809 -604 843 -588
rect 927 588 961 604
rect 927 -604 961 -588
rect 1045 588 1079 604
rect 1045 -604 1079 -588
rect 1163 588 1197 604
rect 1163 -604 1197 -588
rect 1281 588 1315 604
rect 1281 -604 1315 -588
rect 1399 588 1433 604
rect 1399 -604 1433 -588
rect 1517 588 1551 604
rect 1517 -604 1551 -588
rect 1635 588 1669 604
rect 1635 -604 1669 -588
rect 1753 588 1787 604
rect 1753 -604 1787 -588
rect 1871 588 1905 604
rect 1871 -604 1905 -588
rect 1989 588 2023 604
rect 1989 -604 2023 -588
rect 2107 588 2141 604
rect 2107 -604 2141 -588
rect 2225 588 2259 604
rect 2225 -604 2259 -588
rect 2343 588 2377 604
rect 2343 -604 2377 -588
rect 2461 588 2495 604
rect 2461 -604 2495 -588
rect 2579 588 2613 604
rect 2579 -604 2613 -588
rect 2697 588 2731 604
rect 2697 -604 2731 -588
rect 2815 588 2849 604
rect 2815 -604 2849 -588
rect 2933 588 2967 604
rect 2933 -604 2967 -588
rect 3051 588 3085 604
rect 3051 -604 3085 -588
rect 3169 588 3203 604
rect 3169 -604 3203 -588
rect 3287 588 3321 604
rect 3287 -604 3321 -588
rect 3405 588 3439 604
rect 3405 -604 3439 -588
rect 3523 588 3557 604
rect 3523 -604 3557 -588
rect -3514 -681 -3498 -647
rect -3464 -681 -3448 -647
rect -3396 -681 -3380 -647
rect -3346 -681 -3330 -647
rect -3278 -681 -3262 -647
rect -3228 -681 -3212 -647
rect -3160 -681 -3144 -647
rect -3110 -681 -3094 -647
rect -3042 -681 -3026 -647
rect -2992 -681 -2976 -647
rect -2924 -681 -2908 -647
rect -2874 -681 -2858 -647
rect -2806 -681 -2790 -647
rect -2756 -681 -2740 -647
rect -2688 -681 -2672 -647
rect -2638 -681 -2622 -647
rect -2570 -681 -2554 -647
rect -2520 -681 -2504 -647
rect -2452 -681 -2436 -647
rect -2402 -681 -2386 -647
rect -2334 -681 -2318 -647
rect -2284 -681 -2268 -647
rect -2216 -681 -2200 -647
rect -2166 -681 -2150 -647
rect -2098 -681 -2082 -647
rect -2048 -681 -2032 -647
rect -1980 -681 -1964 -647
rect -1930 -681 -1914 -647
rect -1862 -681 -1846 -647
rect -1812 -681 -1796 -647
rect -1744 -681 -1728 -647
rect -1694 -681 -1678 -647
rect -1626 -681 -1610 -647
rect -1576 -681 -1560 -647
rect -1508 -681 -1492 -647
rect -1458 -681 -1442 -647
rect -1390 -681 -1374 -647
rect -1340 -681 -1324 -647
rect -1272 -681 -1256 -647
rect -1222 -681 -1206 -647
rect -1154 -681 -1138 -647
rect -1104 -681 -1088 -647
rect -1036 -681 -1020 -647
rect -986 -681 -970 -647
rect -918 -681 -902 -647
rect -868 -681 -852 -647
rect -800 -681 -784 -647
rect -750 -681 -734 -647
rect -682 -681 -666 -647
rect -632 -681 -616 -647
rect -564 -681 -548 -647
rect -514 -681 -498 -647
rect -446 -681 -430 -647
rect -396 -681 -380 -647
rect -328 -681 -312 -647
rect -278 -681 -262 -647
rect -210 -681 -194 -647
rect -160 -681 -144 -647
rect -92 -681 -76 -647
rect -42 -681 -26 -647
rect 26 -681 42 -647
rect 76 -681 92 -647
rect 144 -681 160 -647
rect 194 -681 210 -647
rect 262 -681 278 -647
rect 312 -681 328 -647
rect 380 -681 396 -647
rect 430 -681 446 -647
rect 498 -681 514 -647
rect 548 -681 564 -647
rect 616 -681 632 -647
rect 666 -681 682 -647
rect 734 -681 750 -647
rect 784 -681 800 -647
rect 852 -681 868 -647
rect 902 -681 918 -647
rect 970 -681 986 -647
rect 1020 -681 1036 -647
rect 1088 -681 1104 -647
rect 1138 -681 1154 -647
rect 1206 -681 1222 -647
rect 1256 -681 1272 -647
rect 1324 -681 1340 -647
rect 1374 -681 1390 -647
rect 1442 -681 1458 -647
rect 1492 -681 1508 -647
rect 1560 -681 1576 -647
rect 1610 -681 1626 -647
rect 1678 -681 1694 -647
rect 1728 -681 1744 -647
rect 1796 -681 1812 -647
rect 1846 -681 1862 -647
rect 1914 -681 1930 -647
rect 1964 -681 1980 -647
rect 2032 -681 2048 -647
rect 2082 -681 2098 -647
rect 2150 -681 2166 -647
rect 2200 -681 2216 -647
rect 2268 -681 2284 -647
rect 2318 -681 2334 -647
rect 2386 -681 2402 -647
rect 2436 -681 2452 -647
rect 2504 -681 2520 -647
rect 2554 -681 2570 -647
rect 2622 -681 2638 -647
rect 2672 -681 2688 -647
rect 2740 -681 2756 -647
rect 2790 -681 2806 -647
rect 2858 -681 2874 -647
rect 2908 -681 2924 -647
rect 2976 -681 2992 -647
rect 3026 -681 3042 -647
rect 3094 -681 3110 -647
rect 3144 -681 3160 -647
rect 3212 -681 3228 -647
rect 3262 -681 3278 -647
rect 3330 -681 3346 -647
rect 3380 -681 3396 -647
rect 3448 -681 3464 -647
rect 3498 -681 3514 -647
<< viali >>
rect -3498 647 -3464 681
rect -3380 647 -3346 681
rect -3262 647 -3228 681
rect -3144 647 -3110 681
rect -3026 647 -2992 681
rect -2908 647 -2874 681
rect -2790 647 -2756 681
rect -2672 647 -2638 681
rect -2554 647 -2520 681
rect -2436 647 -2402 681
rect -2318 647 -2284 681
rect -2200 647 -2166 681
rect -2082 647 -2048 681
rect -1964 647 -1930 681
rect -1846 647 -1812 681
rect -1728 647 -1694 681
rect -1610 647 -1576 681
rect -1492 647 -1458 681
rect -1374 647 -1340 681
rect -1256 647 -1222 681
rect -1138 647 -1104 681
rect -1020 647 -986 681
rect -902 647 -868 681
rect -784 647 -750 681
rect -666 647 -632 681
rect -548 647 -514 681
rect -430 647 -396 681
rect -312 647 -278 681
rect -194 647 -160 681
rect -76 647 -42 681
rect 42 647 76 681
rect 160 647 194 681
rect 278 647 312 681
rect 396 647 430 681
rect 514 647 548 681
rect 632 647 666 681
rect 750 647 784 681
rect 868 647 902 681
rect 986 647 1020 681
rect 1104 647 1138 681
rect 1222 647 1256 681
rect 1340 647 1374 681
rect 1458 647 1492 681
rect 1576 647 1610 681
rect 1694 647 1728 681
rect 1812 647 1846 681
rect 1930 647 1964 681
rect 2048 647 2082 681
rect 2166 647 2200 681
rect 2284 647 2318 681
rect 2402 647 2436 681
rect 2520 647 2554 681
rect 2638 647 2672 681
rect 2756 647 2790 681
rect 2874 647 2908 681
rect 2992 647 3026 681
rect 3110 647 3144 681
rect 3228 647 3262 681
rect 3346 647 3380 681
rect 3464 647 3498 681
rect -3557 -588 -3523 588
rect -3439 -588 -3405 588
rect -3321 -588 -3287 588
rect -3203 -588 -3169 588
rect -3085 -588 -3051 588
rect -2967 -588 -2933 588
rect -2849 -588 -2815 588
rect -2731 -588 -2697 588
rect -2613 -588 -2579 588
rect -2495 -588 -2461 588
rect -2377 -588 -2343 588
rect -2259 -588 -2225 588
rect -2141 -588 -2107 588
rect -2023 -588 -1989 588
rect -1905 -588 -1871 588
rect -1787 -588 -1753 588
rect -1669 -588 -1635 588
rect -1551 -588 -1517 588
rect -1433 -588 -1399 588
rect -1315 -588 -1281 588
rect -1197 -588 -1163 588
rect -1079 -588 -1045 588
rect -961 -588 -927 588
rect -843 -588 -809 588
rect -725 -588 -691 588
rect -607 -588 -573 588
rect -489 -588 -455 588
rect -371 -588 -337 588
rect -253 -588 -219 588
rect -135 -588 -101 588
rect -17 -588 17 588
rect 101 -588 135 588
rect 219 -588 253 588
rect 337 -588 371 588
rect 455 -588 489 588
rect 573 -588 607 588
rect 691 -588 725 588
rect 809 -588 843 588
rect 927 -588 961 588
rect 1045 -588 1079 588
rect 1163 -588 1197 588
rect 1281 -588 1315 588
rect 1399 -588 1433 588
rect 1517 -588 1551 588
rect 1635 -588 1669 588
rect 1753 -588 1787 588
rect 1871 -588 1905 588
rect 1989 -588 2023 588
rect 2107 -588 2141 588
rect 2225 -588 2259 588
rect 2343 -588 2377 588
rect 2461 -588 2495 588
rect 2579 -588 2613 588
rect 2697 -588 2731 588
rect 2815 -588 2849 588
rect 2933 -588 2967 588
rect 3051 -588 3085 588
rect 3169 -588 3203 588
rect 3287 -588 3321 588
rect 3405 -588 3439 588
rect 3523 -588 3557 588
rect -3498 -681 -3464 -647
rect -3380 -681 -3346 -647
rect -3262 -681 -3228 -647
rect -3144 -681 -3110 -647
rect -3026 -681 -2992 -647
rect -2908 -681 -2874 -647
rect -2790 -681 -2756 -647
rect -2672 -681 -2638 -647
rect -2554 -681 -2520 -647
rect -2436 -681 -2402 -647
rect -2318 -681 -2284 -647
rect -2200 -681 -2166 -647
rect -2082 -681 -2048 -647
rect -1964 -681 -1930 -647
rect -1846 -681 -1812 -647
rect -1728 -681 -1694 -647
rect -1610 -681 -1576 -647
rect -1492 -681 -1458 -647
rect -1374 -681 -1340 -647
rect -1256 -681 -1222 -647
rect -1138 -681 -1104 -647
rect -1020 -681 -986 -647
rect -902 -681 -868 -647
rect -784 -681 -750 -647
rect -666 -681 -632 -647
rect -548 -681 -514 -647
rect -430 -681 -396 -647
rect -312 -681 -278 -647
rect -194 -681 -160 -647
rect -76 -681 -42 -647
rect 42 -681 76 -647
rect 160 -681 194 -647
rect 278 -681 312 -647
rect 396 -681 430 -647
rect 514 -681 548 -647
rect 632 -681 666 -647
rect 750 -681 784 -647
rect 868 -681 902 -647
rect 986 -681 1020 -647
rect 1104 -681 1138 -647
rect 1222 -681 1256 -647
rect 1340 -681 1374 -647
rect 1458 -681 1492 -647
rect 1576 -681 1610 -647
rect 1694 -681 1728 -647
rect 1812 -681 1846 -647
rect 1930 -681 1964 -647
rect 2048 -681 2082 -647
rect 2166 -681 2200 -647
rect 2284 -681 2318 -647
rect 2402 -681 2436 -647
rect 2520 -681 2554 -647
rect 2638 -681 2672 -647
rect 2756 -681 2790 -647
rect 2874 -681 2908 -647
rect 2992 -681 3026 -647
rect 3110 -681 3144 -647
rect 3228 -681 3262 -647
rect 3346 -681 3380 -647
rect 3464 -681 3498 -647
<< metal1 >>
rect -3510 681 -3452 687
rect -3510 647 -3498 681
rect -3464 647 -3452 681
rect -3510 641 -3452 647
rect -3392 681 -3334 687
rect -3392 647 -3380 681
rect -3346 647 -3334 681
rect -3392 641 -3334 647
rect -3274 681 -3216 687
rect -3274 647 -3262 681
rect -3228 647 -3216 681
rect -3274 641 -3216 647
rect -3156 681 -3098 687
rect -3156 647 -3144 681
rect -3110 647 -3098 681
rect -3156 641 -3098 647
rect -3038 681 -2980 687
rect -3038 647 -3026 681
rect -2992 647 -2980 681
rect -3038 641 -2980 647
rect -2920 681 -2862 687
rect -2920 647 -2908 681
rect -2874 647 -2862 681
rect -2920 641 -2862 647
rect -2802 681 -2744 687
rect -2802 647 -2790 681
rect -2756 647 -2744 681
rect -2802 641 -2744 647
rect -2684 681 -2626 687
rect -2684 647 -2672 681
rect -2638 647 -2626 681
rect -2684 641 -2626 647
rect -2566 681 -2508 687
rect -2566 647 -2554 681
rect -2520 647 -2508 681
rect -2566 641 -2508 647
rect -2448 681 -2390 687
rect -2448 647 -2436 681
rect -2402 647 -2390 681
rect -2448 641 -2390 647
rect -2330 681 -2272 687
rect -2330 647 -2318 681
rect -2284 647 -2272 681
rect -2330 641 -2272 647
rect -2212 681 -2154 687
rect -2212 647 -2200 681
rect -2166 647 -2154 681
rect -2212 641 -2154 647
rect -2094 681 -2036 687
rect -2094 647 -2082 681
rect -2048 647 -2036 681
rect -2094 641 -2036 647
rect -1976 681 -1918 687
rect -1976 647 -1964 681
rect -1930 647 -1918 681
rect -1976 641 -1918 647
rect -1858 681 -1800 687
rect -1858 647 -1846 681
rect -1812 647 -1800 681
rect -1858 641 -1800 647
rect -1740 681 -1682 687
rect -1740 647 -1728 681
rect -1694 647 -1682 681
rect -1740 641 -1682 647
rect -1622 681 -1564 687
rect -1622 647 -1610 681
rect -1576 647 -1564 681
rect -1622 641 -1564 647
rect -1504 681 -1446 687
rect -1504 647 -1492 681
rect -1458 647 -1446 681
rect -1504 641 -1446 647
rect -1386 681 -1328 687
rect -1386 647 -1374 681
rect -1340 647 -1328 681
rect -1386 641 -1328 647
rect -1268 681 -1210 687
rect -1268 647 -1256 681
rect -1222 647 -1210 681
rect -1268 641 -1210 647
rect -1150 681 -1092 687
rect -1150 647 -1138 681
rect -1104 647 -1092 681
rect -1150 641 -1092 647
rect -1032 681 -974 687
rect -1032 647 -1020 681
rect -986 647 -974 681
rect -1032 641 -974 647
rect -914 681 -856 687
rect -914 647 -902 681
rect -868 647 -856 681
rect -914 641 -856 647
rect -796 681 -738 687
rect -796 647 -784 681
rect -750 647 -738 681
rect -796 641 -738 647
rect -678 681 -620 687
rect -678 647 -666 681
rect -632 647 -620 681
rect -678 641 -620 647
rect -560 681 -502 687
rect -560 647 -548 681
rect -514 647 -502 681
rect -560 641 -502 647
rect -442 681 -384 687
rect -442 647 -430 681
rect -396 647 -384 681
rect -442 641 -384 647
rect -324 681 -266 687
rect -324 647 -312 681
rect -278 647 -266 681
rect -324 641 -266 647
rect -206 681 -148 687
rect -206 647 -194 681
rect -160 647 -148 681
rect -206 641 -148 647
rect -88 681 -30 687
rect -88 647 -76 681
rect -42 647 -30 681
rect -88 641 -30 647
rect 30 681 88 687
rect 30 647 42 681
rect 76 647 88 681
rect 30 641 88 647
rect 148 681 206 687
rect 148 647 160 681
rect 194 647 206 681
rect 148 641 206 647
rect 266 681 324 687
rect 266 647 278 681
rect 312 647 324 681
rect 266 641 324 647
rect 384 681 442 687
rect 384 647 396 681
rect 430 647 442 681
rect 384 641 442 647
rect 502 681 560 687
rect 502 647 514 681
rect 548 647 560 681
rect 502 641 560 647
rect 620 681 678 687
rect 620 647 632 681
rect 666 647 678 681
rect 620 641 678 647
rect 738 681 796 687
rect 738 647 750 681
rect 784 647 796 681
rect 738 641 796 647
rect 856 681 914 687
rect 856 647 868 681
rect 902 647 914 681
rect 856 641 914 647
rect 974 681 1032 687
rect 974 647 986 681
rect 1020 647 1032 681
rect 974 641 1032 647
rect 1092 681 1150 687
rect 1092 647 1104 681
rect 1138 647 1150 681
rect 1092 641 1150 647
rect 1210 681 1268 687
rect 1210 647 1222 681
rect 1256 647 1268 681
rect 1210 641 1268 647
rect 1328 681 1386 687
rect 1328 647 1340 681
rect 1374 647 1386 681
rect 1328 641 1386 647
rect 1446 681 1504 687
rect 1446 647 1458 681
rect 1492 647 1504 681
rect 1446 641 1504 647
rect 1564 681 1622 687
rect 1564 647 1576 681
rect 1610 647 1622 681
rect 1564 641 1622 647
rect 1682 681 1740 687
rect 1682 647 1694 681
rect 1728 647 1740 681
rect 1682 641 1740 647
rect 1800 681 1858 687
rect 1800 647 1812 681
rect 1846 647 1858 681
rect 1800 641 1858 647
rect 1918 681 1976 687
rect 1918 647 1930 681
rect 1964 647 1976 681
rect 1918 641 1976 647
rect 2036 681 2094 687
rect 2036 647 2048 681
rect 2082 647 2094 681
rect 2036 641 2094 647
rect 2154 681 2212 687
rect 2154 647 2166 681
rect 2200 647 2212 681
rect 2154 641 2212 647
rect 2272 681 2330 687
rect 2272 647 2284 681
rect 2318 647 2330 681
rect 2272 641 2330 647
rect 2390 681 2448 687
rect 2390 647 2402 681
rect 2436 647 2448 681
rect 2390 641 2448 647
rect 2508 681 2566 687
rect 2508 647 2520 681
rect 2554 647 2566 681
rect 2508 641 2566 647
rect 2626 681 2684 687
rect 2626 647 2638 681
rect 2672 647 2684 681
rect 2626 641 2684 647
rect 2744 681 2802 687
rect 2744 647 2756 681
rect 2790 647 2802 681
rect 2744 641 2802 647
rect 2862 681 2920 687
rect 2862 647 2874 681
rect 2908 647 2920 681
rect 2862 641 2920 647
rect 2980 681 3038 687
rect 2980 647 2992 681
rect 3026 647 3038 681
rect 2980 641 3038 647
rect 3098 681 3156 687
rect 3098 647 3110 681
rect 3144 647 3156 681
rect 3098 641 3156 647
rect 3216 681 3274 687
rect 3216 647 3228 681
rect 3262 647 3274 681
rect 3216 641 3274 647
rect 3334 681 3392 687
rect 3334 647 3346 681
rect 3380 647 3392 681
rect 3334 641 3392 647
rect 3452 681 3510 687
rect 3452 647 3464 681
rect 3498 647 3510 681
rect 3452 641 3510 647
rect -3563 588 -3517 600
rect -3563 -588 -3557 588
rect -3523 -588 -3517 588
rect -3563 -600 -3517 -588
rect -3445 588 -3399 600
rect -3445 -588 -3439 588
rect -3405 -588 -3399 588
rect -3445 -600 -3399 -588
rect -3327 588 -3281 600
rect -3327 -588 -3321 588
rect -3287 -588 -3281 588
rect -3327 -600 -3281 -588
rect -3209 588 -3163 600
rect -3209 -588 -3203 588
rect -3169 -588 -3163 588
rect -3209 -600 -3163 -588
rect -3091 588 -3045 600
rect -3091 -588 -3085 588
rect -3051 -588 -3045 588
rect -3091 -600 -3045 -588
rect -2973 588 -2927 600
rect -2973 -588 -2967 588
rect -2933 -588 -2927 588
rect -2973 -600 -2927 -588
rect -2855 588 -2809 600
rect -2855 -588 -2849 588
rect -2815 -588 -2809 588
rect -2855 -600 -2809 -588
rect -2737 588 -2691 600
rect -2737 -588 -2731 588
rect -2697 -588 -2691 588
rect -2737 -600 -2691 -588
rect -2619 588 -2573 600
rect -2619 -588 -2613 588
rect -2579 -588 -2573 588
rect -2619 -600 -2573 -588
rect -2501 588 -2455 600
rect -2501 -588 -2495 588
rect -2461 -588 -2455 588
rect -2501 -600 -2455 -588
rect -2383 588 -2337 600
rect -2383 -588 -2377 588
rect -2343 -588 -2337 588
rect -2383 -600 -2337 -588
rect -2265 588 -2219 600
rect -2265 -588 -2259 588
rect -2225 -588 -2219 588
rect -2265 -600 -2219 -588
rect -2147 588 -2101 600
rect -2147 -588 -2141 588
rect -2107 -588 -2101 588
rect -2147 -600 -2101 -588
rect -2029 588 -1983 600
rect -2029 -588 -2023 588
rect -1989 -588 -1983 588
rect -2029 -600 -1983 -588
rect -1911 588 -1865 600
rect -1911 -588 -1905 588
rect -1871 -588 -1865 588
rect -1911 -600 -1865 -588
rect -1793 588 -1747 600
rect -1793 -588 -1787 588
rect -1753 -588 -1747 588
rect -1793 -600 -1747 -588
rect -1675 588 -1629 600
rect -1675 -588 -1669 588
rect -1635 -588 -1629 588
rect -1675 -600 -1629 -588
rect -1557 588 -1511 600
rect -1557 -588 -1551 588
rect -1517 -588 -1511 588
rect -1557 -600 -1511 -588
rect -1439 588 -1393 600
rect -1439 -588 -1433 588
rect -1399 -588 -1393 588
rect -1439 -600 -1393 -588
rect -1321 588 -1275 600
rect -1321 -588 -1315 588
rect -1281 -588 -1275 588
rect -1321 -600 -1275 -588
rect -1203 588 -1157 600
rect -1203 -588 -1197 588
rect -1163 -588 -1157 588
rect -1203 -600 -1157 -588
rect -1085 588 -1039 600
rect -1085 -588 -1079 588
rect -1045 -588 -1039 588
rect -1085 -600 -1039 -588
rect -967 588 -921 600
rect -967 -588 -961 588
rect -927 -588 -921 588
rect -967 -600 -921 -588
rect -849 588 -803 600
rect -849 -588 -843 588
rect -809 -588 -803 588
rect -849 -600 -803 -588
rect -731 588 -685 600
rect -731 -588 -725 588
rect -691 -588 -685 588
rect -731 -600 -685 -588
rect -613 588 -567 600
rect -613 -588 -607 588
rect -573 -588 -567 588
rect -613 -600 -567 -588
rect -495 588 -449 600
rect -495 -588 -489 588
rect -455 -588 -449 588
rect -495 -600 -449 -588
rect -377 588 -331 600
rect -377 -588 -371 588
rect -337 -588 -331 588
rect -377 -600 -331 -588
rect -259 588 -213 600
rect -259 -588 -253 588
rect -219 -588 -213 588
rect -259 -600 -213 -588
rect -141 588 -95 600
rect -141 -588 -135 588
rect -101 -588 -95 588
rect -141 -600 -95 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 95 588 141 600
rect 95 -588 101 588
rect 135 -588 141 588
rect 95 -600 141 -588
rect 213 588 259 600
rect 213 -588 219 588
rect 253 -588 259 588
rect 213 -600 259 -588
rect 331 588 377 600
rect 331 -588 337 588
rect 371 -588 377 588
rect 331 -600 377 -588
rect 449 588 495 600
rect 449 -588 455 588
rect 489 -588 495 588
rect 449 -600 495 -588
rect 567 588 613 600
rect 567 -588 573 588
rect 607 -588 613 588
rect 567 -600 613 -588
rect 685 588 731 600
rect 685 -588 691 588
rect 725 -588 731 588
rect 685 -600 731 -588
rect 803 588 849 600
rect 803 -588 809 588
rect 843 -588 849 588
rect 803 -600 849 -588
rect 921 588 967 600
rect 921 -588 927 588
rect 961 -588 967 588
rect 921 -600 967 -588
rect 1039 588 1085 600
rect 1039 -588 1045 588
rect 1079 -588 1085 588
rect 1039 -600 1085 -588
rect 1157 588 1203 600
rect 1157 -588 1163 588
rect 1197 -588 1203 588
rect 1157 -600 1203 -588
rect 1275 588 1321 600
rect 1275 -588 1281 588
rect 1315 -588 1321 588
rect 1275 -600 1321 -588
rect 1393 588 1439 600
rect 1393 -588 1399 588
rect 1433 -588 1439 588
rect 1393 -600 1439 -588
rect 1511 588 1557 600
rect 1511 -588 1517 588
rect 1551 -588 1557 588
rect 1511 -600 1557 -588
rect 1629 588 1675 600
rect 1629 -588 1635 588
rect 1669 -588 1675 588
rect 1629 -600 1675 -588
rect 1747 588 1793 600
rect 1747 -588 1753 588
rect 1787 -588 1793 588
rect 1747 -600 1793 -588
rect 1865 588 1911 600
rect 1865 -588 1871 588
rect 1905 -588 1911 588
rect 1865 -600 1911 -588
rect 1983 588 2029 600
rect 1983 -588 1989 588
rect 2023 -588 2029 588
rect 1983 -600 2029 -588
rect 2101 588 2147 600
rect 2101 -588 2107 588
rect 2141 -588 2147 588
rect 2101 -600 2147 -588
rect 2219 588 2265 600
rect 2219 -588 2225 588
rect 2259 -588 2265 588
rect 2219 -600 2265 -588
rect 2337 588 2383 600
rect 2337 -588 2343 588
rect 2377 -588 2383 588
rect 2337 -600 2383 -588
rect 2455 588 2501 600
rect 2455 -588 2461 588
rect 2495 -588 2501 588
rect 2455 -600 2501 -588
rect 2573 588 2619 600
rect 2573 -588 2579 588
rect 2613 -588 2619 588
rect 2573 -600 2619 -588
rect 2691 588 2737 600
rect 2691 -588 2697 588
rect 2731 -588 2737 588
rect 2691 -600 2737 -588
rect 2809 588 2855 600
rect 2809 -588 2815 588
rect 2849 -588 2855 588
rect 2809 -600 2855 -588
rect 2927 588 2973 600
rect 2927 -588 2933 588
rect 2967 -588 2973 588
rect 2927 -600 2973 -588
rect 3045 588 3091 600
rect 3045 -588 3051 588
rect 3085 -588 3091 588
rect 3045 -600 3091 -588
rect 3163 588 3209 600
rect 3163 -588 3169 588
rect 3203 -588 3209 588
rect 3163 -600 3209 -588
rect 3281 588 3327 600
rect 3281 -588 3287 588
rect 3321 -588 3327 588
rect 3281 -600 3327 -588
rect 3399 588 3445 600
rect 3399 -588 3405 588
rect 3439 -588 3445 588
rect 3399 -600 3445 -588
rect 3517 588 3563 600
rect 3517 -588 3523 588
rect 3557 -588 3563 588
rect 3517 -600 3563 -588
rect -3510 -647 -3452 -641
rect -3510 -681 -3498 -647
rect -3464 -681 -3452 -647
rect -3510 -687 -3452 -681
rect -3392 -647 -3334 -641
rect -3392 -681 -3380 -647
rect -3346 -681 -3334 -647
rect -3392 -687 -3334 -681
rect -3274 -647 -3216 -641
rect -3274 -681 -3262 -647
rect -3228 -681 -3216 -647
rect -3274 -687 -3216 -681
rect -3156 -647 -3098 -641
rect -3156 -681 -3144 -647
rect -3110 -681 -3098 -647
rect -3156 -687 -3098 -681
rect -3038 -647 -2980 -641
rect -3038 -681 -3026 -647
rect -2992 -681 -2980 -647
rect -3038 -687 -2980 -681
rect -2920 -647 -2862 -641
rect -2920 -681 -2908 -647
rect -2874 -681 -2862 -647
rect -2920 -687 -2862 -681
rect -2802 -647 -2744 -641
rect -2802 -681 -2790 -647
rect -2756 -681 -2744 -647
rect -2802 -687 -2744 -681
rect -2684 -647 -2626 -641
rect -2684 -681 -2672 -647
rect -2638 -681 -2626 -647
rect -2684 -687 -2626 -681
rect -2566 -647 -2508 -641
rect -2566 -681 -2554 -647
rect -2520 -681 -2508 -647
rect -2566 -687 -2508 -681
rect -2448 -647 -2390 -641
rect -2448 -681 -2436 -647
rect -2402 -681 -2390 -647
rect -2448 -687 -2390 -681
rect -2330 -647 -2272 -641
rect -2330 -681 -2318 -647
rect -2284 -681 -2272 -647
rect -2330 -687 -2272 -681
rect -2212 -647 -2154 -641
rect -2212 -681 -2200 -647
rect -2166 -681 -2154 -647
rect -2212 -687 -2154 -681
rect -2094 -647 -2036 -641
rect -2094 -681 -2082 -647
rect -2048 -681 -2036 -647
rect -2094 -687 -2036 -681
rect -1976 -647 -1918 -641
rect -1976 -681 -1964 -647
rect -1930 -681 -1918 -647
rect -1976 -687 -1918 -681
rect -1858 -647 -1800 -641
rect -1858 -681 -1846 -647
rect -1812 -681 -1800 -647
rect -1858 -687 -1800 -681
rect -1740 -647 -1682 -641
rect -1740 -681 -1728 -647
rect -1694 -681 -1682 -647
rect -1740 -687 -1682 -681
rect -1622 -647 -1564 -641
rect -1622 -681 -1610 -647
rect -1576 -681 -1564 -647
rect -1622 -687 -1564 -681
rect -1504 -647 -1446 -641
rect -1504 -681 -1492 -647
rect -1458 -681 -1446 -647
rect -1504 -687 -1446 -681
rect -1386 -647 -1328 -641
rect -1386 -681 -1374 -647
rect -1340 -681 -1328 -647
rect -1386 -687 -1328 -681
rect -1268 -647 -1210 -641
rect -1268 -681 -1256 -647
rect -1222 -681 -1210 -647
rect -1268 -687 -1210 -681
rect -1150 -647 -1092 -641
rect -1150 -681 -1138 -647
rect -1104 -681 -1092 -647
rect -1150 -687 -1092 -681
rect -1032 -647 -974 -641
rect -1032 -681 -1020 -647
rect -986 -681 -974 -647
rect -1032 -687 -974 -681
rect -914 -647 -856 -641
rect -914 -681 -902 -647
rect -868 -681 -856 -647
rect -914 -687 -856 -681
rect -796 -647 -738 -641
rect -796 -681 -784 -647
rect -750 -681 -738 -647
rect -796 -687 -738 -681
rect -678 -647 -620 -641
rect -678 -681 -666 -647
rect -632 -681 -620 -647
rect -678 -687 -620 -681
rect -560 -647 -502 -641
rect -560 -681 -548 -647
rect -514 -681 -502 -647
rect -560 -687 -502 -681
rect -442 -647 -384 -641
rect -442 -681 -430 -647
rect -396 -681 -384 -647
rect -442 -687 -384 -681
rect -324 -647 -266 -641
rect -324 -681 -312 -647
rect -278 -681 -266 -647
rect -324 -687 -266 -681
rect -206 -647 -148 -641
rect -206 -681 -194 -647
rect -160 -681 -148 -647
rect -206 -687 -148 -681
rect -88 -647 -30 -641
rect -88 -681 -76 -647
rect -42 -681 -30 -647
rect -88 -687 -30 -681
rect 30 -647 88 -641
rect 30 -681 42 -647
rect 76 -681 88 -647
rect 30 -687 88 -681
rect 148 -647 206 -641
rect 148 -681 160 -647
rect 194 -681 206 -647
rect 148 -687 206 -681
rect 266 -647 324 -641
rect 266 -681 278 -647
rect 312 -681 324 -647
rect 266 -687 324 -681
rect 384 -647 442 -641
rect 384 -681 396 -647
rect 430 -681 442 -647
rect 384 -687 442 -681
rect 502 -647 560 -641
rect 502 -681 514 -647
rect 548 -681 560 -647
rect 502 -687 560 -681
rect 620 -647 678 -641
rect 620 -681 632 -647
rect 666 -681 678 -647
rect 620 -687 678 -681
rect 738 -647 796 -641
rect 738 -681 750 -647
rect 784 -681 796 -647
rect 738 -687 796 -681
rect 856 -647 914 -641
rect 856 -681 868 -647
rect 902 -681 914 -647
rect 856 -687 914 -681
rect 974 -647 1032 -641
rect 974 -681 986 -647
rect 1020 -681 1032 -647
rect 974 -687 1032 -681
rect 1092 -647 1150 -641
rect 1092 -681 1104 -647
rect 1138 -681 1150 -647
rect 1092 -687 1150 -681
rect 1210 -647 1268 -641
rect 1210 -681 1222 -647
rect 1256 -681 1268 -647
rect 1210 -687 1268 -681
rect 1328 -647 1386 -641
rect 1328 -681 1340 -647
rect 1374 -681 1386 -647
rect 1328 -687 1386 -681
rect 1446 -647 1504 -641
rect 1446 -681 1458 -647
rect 1492 -681 1504 -647
rect 1446 -687 1504 -681
rect 1564 -647 1622 -641
rect 1564 -681 1576 -647
rect 1610 -681 1622 -647
rect 1564 -687 1622 -681
rect 1682 -647 1740 -641
rect 1682 -681 1694 -647
rect 1728 -681 1740 -647
rect 1682 -687 1740 -681
rect 1800 -647 1858 -641
rect 1800 -681 1812 -647
rect 1846 -681 1858 -647
rect 1800 -687 1858 -681
rect 1918 -647 1976 -641
rect 1918 -681 1930 -647
rect 1964 -681 1976 -647
rect 1918 -687 1976 -681
rect 2036 -647 2094 -641
rect 2036 -681 2048 -647
rect 2082 -681 2094 -647
rect 2036 -687 2094 -681
rect 2154 -647 2212 -641
rect 2154 -681 2166 -647
rect 2200 -681 2212 -647
rect 2154 -687 2212 -681
rect 2272 -647 2330 -641
rect 2272 -681 2284 -647
rect 2318 -681 2330 -647
rect 2272 -687 2330 -681
rect 2390 -647 2448 -641
rect 2390 -681 2402 -647
rect 2436 -681 2448 -647
rect 2390 -687 2448 -681
rect 2508 -647 2566 -641
rect 2508 -681 2520 -647
rect 2554 -681 2566 -647
rect 2508 -687 2566 -681
rect 2626 -647 2684 -641
rect 2626 -681 2638 -647
rect 2672 -681 2684 -647
rect 2626 -687 2684 -681
rect 2744 -647 2802 -641
rect 2744 -681 2756 -647
rect 2790 -681 2802 -647
rect 2744 -687 2802 -681
rect 2862 -647 2920 -641
rect 2862 -681 2874 -647
rect 2908 -681 2920 -647
rect 2862 -687 2920 -681
rect 2980 -647 3038 -641
rect 2980 -681 2992 -647
rect 3026 -681 3038 -647
rect 2980 -687 3038 -681
rect 3098 -647 3156 -641
rect 3098 -681 3110 -647
rect 3144 -681 3156 -647
rect 3098 -687 3156 -681
rect 3216 -647 3274 -641
rect 3216 -681 3228 -647
rect 3262 -681 3274 -647
rect 3216 -687 3274 -681
rect 3334 -647 3392 -641
rect 3334 -681 3346 -647
rect 3380 -681 3392 -647
rect 3334 -687 3392 -681
rect 3452 -647 3510 -641
rect 3452 -681 3464 -647
rect 3498 -681 3510 -647
rect 3452 -687 3510 -681
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.3 m 1 nf 60 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
