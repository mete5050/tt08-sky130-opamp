magic
tech sky130B
timestamp 1768737176
<< nmos >>
rect -179 -299 -79 268
rect -50 -299 50 268
rect 79 -299 179 268
<< ndiff >>
rect -208 262 -179 268
rect -208 -293 -202 262
rect -185 -293 -179 262
rect -208 -299 -179 -293
rect -79 262 -50 268
rect -79 -293 -73 262
rect -56 -293 -50 262
rect -79 -299 -50 -293
rect 50 262 79 268
rect 50 -293 56 262
rect 73 -293 79 262
rect 50 -299 79 -293
rect 179 262 208 268
rect 179 -293 185 262
rect 202 -293 208 262
rect 179 -299 208 -293
<< ndiffc >>
rect -202 -293 -185 262
rect -73 -293 -56 262
rect 56 -293 73 262
rect 185 -293 202 262
<< poly >>
rect -179 304 -79 312
rect -179 287 -171 304
rect -87 287 -79 304
rect -179 268 -79 287
rect -50 304 50 312
rect -50 287 -42 304
rect 42 287 50 304
rect -50 268 50 287
rect 79 304 179 312
rect 79 287 87 304
rect 171 287 179 304
rect 79 268 179 287
rect -179 -312 -79 -299
rect -50 -312 50 -299
rect 79 -312 179 -299
<< polycont >>
rect -171 287 -87 304
rect -42 287 42 304
rect 87 287 171 304
<< locali >>
rect -179 287 -171 304
rect -87 287 -79 304
rect -50 287 -42 304
rect 42 287 50 304
rect 79 287 87 304
rect 171 287 179 304
rect -202 262 -185 270
rect -202 -301 -185 -293
rect -73 262 -56 270
rect -73 -301 -56 -293
rect 56 262 73 270
rect 56 -301 73 -293
rect 185 262 202 270
rect 185 -301 202 -293
<< viali >>
rect -171 287 -87 304
rect -42 287 42 304
rect 87 287 171 304
rect -202 -293 -185 262
rect -73 -293 -56 262
rect 56 -293 73 262
rect 185 -293 202 262
<< metal1 >>
rect -177 304 -81 307
rect -177 287 -171 304
rect -87 287 -81 304
rect -177 284 -81 287
rect -48 304 48 307
rect -48 287 -42 304
rect 42 287 48 304
rect -48 284 48 287
rect 81 304 177 307
rect 81 287 87 304
rect 171 287 177 304
rect 81 284 177 287
rect -205 262 -182 268
rect -205 -293 -202 262
rect -185 -293 -182 262
rect -205 -299 -182 -293
rect -76 262 -53 268
rect -76 -293 -73 262
rect -56 -293 -53 262
rect -76 -299 -53 -293
rect 53 262 76 268
rect 53 -293 56 262
rect 73 -293 76 262
rect 53 -299 76 -293
rect 182 262 205 268
rect 182 -293 185 262
rect 202 -293 205 262
rect 182 -299 205 -293
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.666666666666667 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
