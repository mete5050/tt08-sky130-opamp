magic
tech sky130B
magscale 1 2
timestamp 1768749944
<< nmos >>
rect -100 -131 100 69
<< ndiff >>
rect -158 57 -100 69
rect -158 -119 -146 57
rect -112 -119 -100 57
rect -158 -131 -100 -119
rect 100 57 158 69
rect 100 -119 112 57
rect 146 -119 158 57
rect 100 -131 158 -119
<< ndiffc >>
rect -146 -119 -112 57
rect 112 -119 146 57
<< poly >>
rect -100 141 100 157
rect -100 107 -84 141
rect 84 107 100 141
rect -100 69 100 107
rect -100 -157 100 -131
<< polycont >>
rect -84 107 84 141
<< locali >>
rect -100 107 -84 141
rect 84 107 100 141
rect -146 57 -112 73
rect -146 -135 -112 -119
rect 112 57 146 73
rect 112 -135 146 -119
<< viali >>
rect -84 107 84 141
rect -146 -119 -112 57
rect 112 -119 146 57
<< metal1 >>
rect -96 141 96 147
rect -96 107 -84 141
rect 84 107 96 141
rect -96 101 96 107
rect -152 57 -106 69
rect -152 -119 -146 57
rect -112 -119 -106 57
rect -152 -131 -106 -119
rect 106 57 152 69
rect 106 -119 112 57
rect 146 -119 152 57
rect 106 -131 152 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
