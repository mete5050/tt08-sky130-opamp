magic
tech sky130B
magscale 1 2
timestamp 1768750829
<< nmos >>
rect -616 -569 -416 631
rect -358 -569 -158 631
rect -100 -569 100 631
rect 158 -569 358 631
rect 416 -569 616 631
<< ndiff >>
rect -674 619 -616 631
rect -674 -557 -662 619
rect -628 -557 -616 619
rect -674 -569 -616 -557
rect -416 619 -358 631
rect -416 -557 -404 619
rect -370 -557 -358 619
rect -416 -569 -358 -557
rect -158 619 -100 631
rect -158 -557 -146 619
rect -112 -557 -100 619
rect -158 -569 -100 -557
rect 100 619 158 631
rect 100 -557 112 619
rect 146 -557 158 619
rect 100 -569 158 -557
rect 358 619 416 631
rect 358 -557 370 619
rect 404 -557 416 619
rect 358 -569 416 -557
rect 616 619 674 631
rect 616 -557 628 619
rect 662 -557 674 619
rect 616 -569 674 -557
<< ndiffc >>
rect -662 -557 -628 619
rect -404 -557 -370 619
rect -146 -557 -112 619
rect 112 -557 146 619
rect 370 -557 404 619
rect 628 -557 662 619
<< poly >>
rect -616 631 -416 657
rect -358 631 -158 657
rect -100 631 100 657
rect 158 631 358 657
rect 416 631 616 657
rect -616 -607 -416 -569
rect -616 -641 -600 -607
rect -432 -641 -416 -607
rect -616 -657 -416 -641
rect -358 -607 -158 -569
rect -358 -641 -342 -607
rect -174 -641 -158 -607
rect -358 -657 -158 -641
rect -100 -607 100 -569
rect -100 -641 -84 -607
rect 84 -641 100 -607
rect -100 -657 100 -641
rect 158 -607 358 -569
rect 158 -641 174 -607
rect 342 -641 358 -607
rect 158 -657 358 -641
rect 416 -607 616 -569
rect 416 -641 432 -607
rect 600 -641 616 -607
rect 416 -657 616 -641
<< polycont >>
rect -600 -641 -432 -607
rect -342 -641 -174 -607
rect -84 -641 84 -607
rect 174 -641 342 -607
rect 432 -641 600 -607
<< locali >>
rect -662 619 -628 635
rect -662 -573 -628 -557
rect -404 619 -370 635
rect -404 -573 -370 -557
rect -146 619 -112 635
rect -146 -573 -112 -557
rect 112 619 146 635
rect 112 -573 146 -557
rect 370 619 404 635
rect 370 -573 404 -557
rect 628 619 662 635
rect 628 -573 662 -557
rect -616 -641 -600 -607
rect -432 -641 -416 -607
rect -358 -641 -342 -607
rect -174 -641 -158 -607
rect -100 -641 -84 -607
rect 84 -641 100 -607
rect 158 -641 174 -607
rect 342 -641 358 -607
rect 416 -641 432 -607
rect 600 -641 616 -607
<< viali >>
rect -662 -557 -628 619
rect -404 -557 -370 619
rect -146 -557 -112 619
rect 112 -557 146 619
rect 370 -557 404 619
rect 628 -557 662 619
rect -600 -641 -432 -607
rect -342 -641 -174 -607
rect -84 -641 84 -607
rect 174 -641 342 -607
rect 432 -641 600 -607
<< metal1 >>
rect -668 619 -622 631
rect -668 -557 -662 619
rect -628 -557 -622 619
rect -668 -569 -622 -557
rect -410 619 -364 631
rect -410 -557 -404 619
rect -370 -557 -364 619
rect -410 -569 -364 -557
rect -152 619 -106 631
rect -152 -557 -146 619
rect -112 -557 -106 619
rect -152 -569 -106 -557
rect 106 619 152 631
rect 106 -557 112 619
rect 146 -557 152 619
rect 106 -569 152 -557
rect 364 619 410 631
rect 364 -557 370 619
rect 404 -557 410 619
rect 364 -569 410 -557
rect 622 619 668 631
rect 622 -557 628 619
rect 662 -557 668 619
rect 622 -569 668 -557
rect -612 -607 -420 -601
rect -612 -641 -600 -607
rect -432 -641 -420 -607
rect -612 -647 -420 -641
rect -354 -607 -162 -601
rect -354 -641 -342 -607
rect -174 -641 -162 -607
rect -354 -647 -162 -641
rect -96 -607 96 -601
rect -96 -641 -84 -607
rect 84 -641 96 -607
rect -96 -647 96 -641
rect 162 -607 354 -601
rect 162 -641 174 -607
rect 342 -641 354 -607
rect 162 -647 354 -641
rect 420 -607 612 -601
rect 420 -641 432 -607
rect 600 -641 612 -607
rect 420 -647 612 -641
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
