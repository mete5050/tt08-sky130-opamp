magic
tech sky130B
magscale 1 2
timestamp 1768734963
<< nwell >>
rect -812 -819 812 819
<< pmos >>
rect -616 -600 -416 600
rect -358 -600 -158 600
rect -100 -600 100 600
rect 158 -600 358 600
rect 416 -600 616 600
<< pdiff >>
rect -674 588 -616 600
rect -674 -588 -662 588
rect -628 -588 -616 588
rect -674 -600 -616 -588
rect -416 588 -358 600
rect -416 -588 -404 588
rect -370 -588 -358 588
rect -416 -600 -358 -588
rect -158 588 -100 600
rect -158 -588 -146 588
rect -112 -588 -100 588
rect -158 -600 -100 -588
rect 100 588 158 600
rect 100 -588 112 588
rect 146 -588 158 588
rect 100 -600 158 -588
rect 358 588 416 600
rect 358 -588 370 588
rect 404 -588 416 588
rect 358 -600 416 -588
rect 616 588 674 600
rect 616 -588 628 588
rect 662 -588 674 588
rect 616 -600 674 -588
<< pdiffc >>
rect -662 -588 -628 588
rect -404 -588 -370 588
rect -146 -588 -112 588
rect 112 -588 146 588
rect 370 -588 404 588
rect 628 -588 662 588
<< nsubdiff >>
rect -776 749 -680 783
rect 680 749 776 783
rect -776 687 -742 749
rect 742 687 776 749
rect -776 -749 -742 -687
rect 742 -749 776 -687
rect -776 -783 -680 -749
rect 680 -783 776 -749
<< nsubdiffcont >>
rect -680 749 680 783
rect -776 -687 -742 687
rect 742 -687 776 687
rect -680 -783 680 -749
<< poly >>
rect -616 681 -416 697
rect -616 647 -600 681
rect -432 647 -416 681
rect -616 600 -416 647
rect -358 681 -158 697
rect -358 647 -342 681
rect -174 647 -158 681
rect -358 600 -158 647
rect -100 681 100 697
rect -100 647 -84 681
rect 84 647 100 681
rect -100 600 100 647
rect 158 681 358 697
rect 158 647 174 681
rect 342 647 358 681
rect 158 600 358 647
rect 416 681 616 697
rect 416 647 432 681
rect 600 647 616 681
rect 416 600 616 647
rect -616 -647 -416 -600
rect -616 -681 -600 -647
rect -432 -681 -416 -647
rect -616 -697 -416 -681
rect -358 -647 -158 -600
rect -358 -681 -342 -647
rect -174 -681 -158 -647
rect -358 -697 -158 -681
rect -100 -647 100 -600
rect -100 -681 -84 -647
rect 84 -681 100 -647
rect -100 -697 100 -681
rect 158 -647 358 -600
rect 158 -681 174 -647
rect 342 -681 358 -647
rect 158 -697 358 -681
rect 416 -647 616 -600
rect 416 -681 432 -647
rect 600 -681 616 -647
rect 416 -697 616 -681
<< polycont >>
rect -600 647 -432 681
rect -342 647 -174 681
rect -84 647 84 681
rect 174 647 342 681
rect 432 647 600 681
rect -600 -681 -432 -647
rect -342 -681 -174 -647
rect -84 -681 84 -647
rect 174 -681 342 -647
rect 432 -681 600 -647
<< locali >>
rect -776 749 -680 783
rect 680 749 776 783
rect -776 687 -742 749
rect 742 687 776 749
rect -616 647 -600 681
rect -432 647 -416 681
rect -358 647 -342 681
rect -174 647 -158 681
rect -100 647 -84 681
rect 84 647 100 681
rect 158 647 174 681
rect 342 647 358 681
rect 416 647 432 681
rect 600 647 616 681
rect -662 588 -628 604
rect -662 -604 -628 -588
rect -404 588 -370 604
rect -404 -604 -370 -588
rect -146 588 -112 604
rect -146 -604 -112 -588
rect 112 588 146 604
rect 112 -604 146 -588
rect 370 588 404 604
rect 370 -604 404 -588
rect 628 588 662 604
rect 628 -604 662 -588
rect -616 -681 -600 -647
rect -432 -681 -416 -647
rect -358 -681 -342 -647
rect -174 -681 -158 -647
rect -100 -681 -84 -647
rect 84 -681 100 -647
rect 158 -681 174 -647
rect 342 -681 358 -647
rect 416 -681 432 -647
rect 600 -681 616 -647
rect -776 -749 -742 -687
rect 742 -749 776 -687
rect -776 -783 -680 -749
rect 680 -783 776 -749
<< viali >>
rect -600 647 -432 681
rect -342 647 -174 681
rect -84 647 84 681
rect 174 647 342 681
rect 432 647 600 681
rect -662 -588 -628 588
rect -404 -588 -370 588
rect -146 -588 -112 588
rect 112 -588 146 588
rect 370 -588 404 588
rect 628 -588 662 588
rect -600 -681 -432 -647
rect -342 -681 -174 -647
rect -84 -681 84 -647
rect 174 -681 342 -647
rect 432 -681 600 -647
<< metal1 >>
rect -612 681 -420 687
rect -612 647 -600 681
rect -432 647 -420 681
rect -612 641 -420 647
rect -354 681 -162 687
rect -354 647 -342 681
rect -174 647 -162 681
rect -354 641 -162 647
rect -96 681 96 687
rect -96 647 -84 681
rect 84 647 96 681
rect -96 641 96 647
rect 162 681 354 687
rect 162 647 174 681
rect 342 647 354 681
rect 162 641 354 647
rect 420 681 612 687
rect 420 647 432 681
rect 600 647 612 681
rect 420 641 612 647
rect -668 588 -622 600
rect -668 -588 -662 588
rect -628 -588 -622 588
rect -668 -600 -622 -588
rect -410 588 -364 600
rect -410 -588 -404 588
rect -370 -588 -364 588
rect -410 -600 -364 -588
rect -152 588 -106 600
rect -152 -588 -146 588
rect -112 -588 -106 588
rect -152 -600 -106 -588
rect 106 588 152 600
rect 106 -588 112 588
rect 146 -588 152 588
rect 106 -600 152 -588
rect 364 588 410 600
rect 364 -588 370 588
rect 404 -588 410 588
rect 364 -600 410 -588
rect 622 588 668 600
rect 622 -588 628 588
rect 662 -588 668 588
rect 622 -600 668 -588
rect -612 -647 -420 -641
rect -612 -681 -600 -647
rect -432 -681 -420 -647
rect -612 -687 -420 -681
rect -354 -647 -162 -641
rect -354 -681 -342 -647
rect -174 -681 -162 -647
rect -354 -687 -162 -681
rect -96 -647 96 -641
rect -96 -681 -84 -647
rect 84 -681 96 -647
rect -96 -687 96 -681
rect 162 -647 354 -641
rect 162 -681 174 -647
rect 342 -681 354 -647
rect 162 -687 354 -681
rect 420 -647 612 -641
rect 420 -681 432 -647
rect 600 -681 612 -647
rect 420 -687 612 -681
<< properties >>
string FIXED_BBOX -759 -766 759 766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
