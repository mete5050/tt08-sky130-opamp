magic
tech sky130B
magscale 1 2
timestamp 1768735973
<< nwell >>
rect -710 -698 710 664
<< pmos >>
rect -616 -636 -416 564
rect -358 -636 -158 564
rect -100 -636 100 564
rect 158 -636 358 564
rect 416 -636 616 564
<< pdiff >>
rect -674 552 -616 564
rect -674 -624 -662 552
rect -628 -624 -616 552
rect -674 -636 -616 -624
rect -416 552 -358 564
rect -416 -624 -404 552
rect -370 -624 -358 552
rect -416 -636 -358 -624
rect -158 552 -100 564
rect -158 -624 -146 552
rect -112 -624 -100 552
rect -158 -636 -100 -624
rect 100 552 158 564
rect 100 -624 112 552
rect 146 -624 158 552
rect 100 -636 158 -624
rect 358 552 416 564
rect 358 -624 370 552
rect 404 -624 416 552
rect 358 -636 416 -624
rect 616 552 674 564
rect 616 -624 628 552
rect 662 -624 674 552
rect 616 -636 674 -624
<< pdiffc >>
rect -662 -624 -628 552
rect -404 -624 -370 552
rect -146 -624 -112 552
rect 112 -624 146 552
rect 370 -624 404 552
rect 628 -624 662 552
<< poly >>
rect -616 645 -416 661
rect -616 611 -600 645
rect -432 611 -416 645
rect -616 564 -416 611
rect -358 645 -158 661
rect -358 611 -342 645
rect -174 611 -158 645
rect -358 564 -158 611
rect -100 645 100 661
rect -100 611 -84 645
rect 84 611 100 645
rect -100 564 100 611
rect 158 645 358 661
rect 158 611 174 645
rect 342 611 358 645
rect 158 564 358 611
rect 416 645 616 661
rect 416 611 432 645
rect 600 611 616 645
rect 416 564 616 611
rect -616 -662 -416 -636
rect -358 -662 -158 -636
rect -100 -662 100 -636
rect 158 -662 358 -636
rect 416 -662 616 -636
<< polycont >>
rect -600 611 -432 645
rect -342 611 -174 645
rect -84 611 84 645
rect 174 611 342 645
rect 432 611 600 645
<< locali >>
rect -616 611 -600 645
rect -432 611 -416 645
rect -358 611 -342 645
rect -174 611 -158 645
rect -100 611 -84 645
rect 84 611 100 645
rect 158 611 174 645
rect 342 611 358 645
rect 416 611 432 645
rect 600 611 616 645
rect -662 552 -628 568
rect -662 -640 -628 -624
rect -404 552 -370 568
rect -404 -640 -370 -624
rect -146 552 -112 568
rect -146 -640 -112 -624
rect 112 552 146 568
rect 112 -640 146 -624
rect 370 552 404 568
rect 370 -640 404 -624
rect 628 552 662 568
rect 628 -640 662 -624
<< viali >>
rect -600 611 -432 645
rect -342 611 -174 645
rect -84 611 84 645
rect 174 611 342 645
rect 432 611 600 645
rect -662 -624 -628 552
rect -404 -624 -370 552
rect -146 -624 -112 552
rect 112 -624 146 552
rect 370 -624 404 552
rect 628 -624 662 552
<< metal1 >>
rect -612 645 -420 651
rect -612 611 -600 645
rect -432 611 -420 645
rect -612 605 -420 611
rect -354 645 -162 651
rect -354 611 -342 645
rect -174 611 -162 645
rect -354 605 -162 611
rect -96 645 96 651
rect -96 611 -84 645
rect 84 611 96 645
rect -96 605 96 611
rect 162 645 354 651
rect 162 611 174 645
rect 342 611 354 645
rect 162 605 354 611
rect 420 645 612 651
rect 420 611 432 645
rect 600 611 612 645
rect 420 605 612 611
rect -668 552 -622 564
rect -668 -624 -662 552
rect -628 -624 -622 552
rect -668 -636 -622 -624
rect -410 552 -364 564
rect -410 -624 -404 552
rect -370 -624 -364 552
rect -410 -636 -364 -624
rect -152 552 -106 564
rect -152 -624 -146 552
rect -112 -624 -106 552
rect -152 -636 -106 -624
rect 106 552 152 564
rect 106 -624 112 552
rect 146 -624 152 552
rect 106 -636 152 -624
rect 364 552 410 564
rect 364 -624 370 552
rect 404 -624 410 552
rect 364 -636 410 -624
rect 622 552 668 564
rect 622 -624 628 552
rect 662 -624 668 552
rect 622 -636 668 -624
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
