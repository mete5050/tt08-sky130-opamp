magic
tech sky130B
magscale 1 2
timestamp 1768735447
<< nwell >>
rect -1355 -664 1355 698
<< pmos >>
rect -1261 -564 -1061 636
rect -1003 -564 -803 636
rect -745 -564 -545 636
rect -487 -564 -287 636
rect -229 -564 -29 636
rect 29 -564 229 636
rect 287 -564 487 636
rect 545 -564 745 636
rect 803 -564 1003 636
rect 1061 -564 1261 636
<< pdiff >>
rect -1319 624 -1261 636
rect -1319 -552 -1307 624
rect -1273 -552 -1261 624
rect -1319 -564 -1261 -552
rect -1061 624 -1003 636
rect -1061 -552 -1049 624
rect -1015 -552 -1003 624
rect -1061 -564 -1003 -552
rect -803 624 -745 636
rect -803 -552 -791 624
rect -757 -552 -745 624
rect -803 -564 -745 -552
rect -545 624 -487 636
rect -545 -552 -533 624
rect -499 -552 -487 624
rect -545 -564 -487 -552
rect -287 624 -229 636
rect -287 -552 -275 624
rect -241 -552 -229 624
rect -287 -564 -229 -552
rect -29 624 29 636
rect -29 -552 -17 624
rect 17 -552 29 624
rect -29 -564 29 -552
rect 229 624 287 636
rect 229 -552 241 624
rect 275 -552 287 624
rect 229 -564 287 -552
rect 487 624 545 636
rect 487 -552 499 624
rect 533 -552 545 624
rect 487 -564 545 -552
rect 745 624 803 636
rect 745 -552 757 624
rect 791 -552 803 624
rect 745 -564 803 -552
rect 1003 624 1061 636
rect 1003 -552 1015 624
rect 1049 -552 1061 624
rect 1003 -564 1061 -552
rect 1261 624 1319 636
rect 1261 -552 1273 624
rect 1307 -552 1319 624
rect 1261 -564 1319 -552
<< pdiffc >>
rect -1307 -552 -1273 624
rect -1049 -552 -1015 624
rect -791 -552 -757 624
rect -533 -552 -499 624
rect -275 -552 -241 624
rect -17 -552 17 624
rect 241 -552 275 624
rect 499 -552 533 624
rect 757 -552 791 624
rect 1015 -552 1049 624
rect 1273 -552 1307 624
<< poly >>
rect -1261 636 -1061 662
rect -1003 636 -803 662
rect -745 636 -545 662
rect -487 636 -287 662
rect -229 636 -29 662
rect 29 636 229 662
rect 287 636 487 662
rect 545 636 745 662
rect 803 636 1003 662
rect 1061 636 1261 662
rect -1261 -611 -1061 -564
rect -1261 -645 -1245 -611
rect -1077 -645 -1061 -611
rect -1261 -661 -1061 -645
rect -1003 -611 -803 -564
rect -1003 -645 -987 -611
rect -819 -645 -803 -611
rect -1003 -661 -803 -645
rect -745 -611 -545 -564
rect -745 -645 -729 -611
rect -561 -645 -545 -611
rect -745 -661 -545 -645
rect -487 -611 -287 -564
rect -487 -645 -471 -611
rect -303 -645 -287 -611
rect -487 -661 -287 -645
rect -229 -611 -29 -564
rect -229 -645 -213 -611
rect -45 -645 -29 -611
rect -229 -661 -29 -645
rect 29 -611 229 -564
rect 29 -645 45 -611
rect 213 -645 229 -611
rect 29 -661 229 -645
rect 287 -611 487 -564
rect 287 -645 303 -611
rect 471 -645 487 -611
rect 287 -661 487 -645
rect 545 -611 745 -564
rect 545 -645 561 -611
rect 729 -645 745 -611
rect 545 -661 745 -645
rect 803 -611 1003 -564
rect 803 -645 819 -611
rect 987 -645 1003 -611
rect 803 -661 1003 -645
rect 1061 -611 1261 -564
rect 1061 -645 1077 -611
rect 1245 -645 1261 -611
rect 1061 -661 1261 -645
<< polycont >>
rect -1245 -645 -1077 -611
rect -987 -645 -819 -611
rect -729 -645 -561 -611
rect -471 -645 -303 -611
rect -213 -645 -45 -611
rect 45 -645 213 -611
rect 303 -645 471 -611
rect 561 -645 729 -611
rect 819 -645 987 -611
rect 1077 -645 1245 -611
<< locali >>
rect -1307 624 -1273 640
rect -1307 -568 -1273 -552
rect -1049 624 -1015 640
rect -1049 -568 -1015 -552
rect -791 624 -757 640
rect -791 -568 -757 -552
rect -533 624 -499 640
rect -533 -568 -499 -552
rect -275 624 -241 640
rect -275 -568 -241 -552
rect -17 624 17 640
rect -17 -568 17 -552
rect 241 624 275 640
rect 241 -568 275 -552
rect 499 624 533 640
rect 499 -568 533 -552
rect 757 624 791 640
rect 757 -568 791 -552
rect 1015 624 1049 640
rect 1015 -568 1049 -552
rect 1273 624 1307 640
rect 1273 -568 1307 -552
rect -1261 -645 -1245 -611
rect -1077 -645 -1061 -611
rect -1003 -645 -987 -611
rect -819 -645 -803 -611
rect -745 -645 -729 -611
rect -561 -645 -545 -611
rect -487 -645 -471 -611
rect -303 -645 -287 -611
rect -229 -645 -213 -611
rect -45 -645 -29 -611
rect 29 -645 45 -611
rect 213 -645 229 -611
rect 287 -645 303 -611
rect 471 -645 487 -611
rect 545 -645 561 -611
rect 729 -645 745 -611
rect 803 -645 819 -611
rect 987 -645 1003 -611
rect 1061 -645 1077 -611
rect 1245 -645 1261 -611
<< viali >>
rect -1307 -552 -1273 624
rect -1049 -552 -1015 624
rect -791 -552 -757 624
rect -533 -552 -499 624
rect -275 -552 -241 624
rect -17 -552 17 624
rect 241 -552 275 624
rect 499 -552 533 624
rect 757 -552 791 624
rect 1015 -552 1049 624
rect 1273 -552 1307 624
rect -1245 -645 -1077 -611
rect -987 -645 -819 -611
rect -729 -645 -561 -611
rect -471 -645 -303 -611
rect -213 -645 -45 -611
rect 45 -645 213 -611
rect 303 -645 471 -611
rect 561 -645 729 -611
rect 819 -645 987 -611
rect 1077 -645 1245 -611
<< metal1 >>
rect -1313 624 -1267 636
rect -1313 -552 -1307 624
rect -1273 -552 -1267 624
rect -1313 -564 -1267 -552
rect -1055 624 -1009 636
rect -1055 -552 -1049 624
rect -1015 -552 -1009 624
rect -1055 -564 -1009 -552
rect -797 624 -751 636
rect -797 -552 -791 624
rect -757 -552 -751 624
rect -797 -564 -751 -552
rect -539 624 -493 636
rect -539 -552 -533 624
rect -499 -552 -493 624
rect -539 -564 -493 -552
rect -281 624 -235 636
rect -281 -552 -275 624
rect -241 -552 -235 624
rect -281 -564 -235 -552
rect -23 624 23 636
rect -23 -552 -17 624
rect 17 -552 23 624
rect -23 -564 23 -552
rect 235 624 281 636
rect 235 -552 241 624
rect 275 -552 281 624
rect 235 -564 281 -552
rect 493 624 539 636
rect 493 -552 499 624
rect 533 -552 539 624
rect 493 -564 539 -552
rect 751 624 797 636
rect 751 -552 757 624
rect 791 -552 797 624
rect 751 -564 797 -552
rect 1009 624 1055 636
rect 1009 -552 1015 624
rect 1049 -552 1055 624
rect 1009 -564 1055 -552
rect 1267 624 1313 636
rect 1267 -552 1273 624
rect 1307 -552 1313 624
rect 1267 -564 1313 -552
rect -1257 -611 -1065 -605
rect -1257 -645 -1245 -611
rect -1077 -645 -1065 -611
rect -1257 -651 -1065 -645
rect -999 -611 -807 -605
rect -999 -645 -987 -611
rect -819 -645 -807 -611
rect -999 -651 -807 -645
rect -741 -611 -549 -605
rect -741 -645 -729 -611
rect -561 -645 -549 -611
rect -741 -651 -549 -645
rect -483 -611 -291 -605
rect -483 -645 -471 -611
rect -303 -645 -291 -611
rect -483 -651 -291 -645
rect -225 -611 -33 -605
rect -225 -645 -213 -611
rect -45 -645 -33 -611
rect -225 -651 -33 -645
rect 33 -611 225 -605
rect 33 -645 45 -611
rect 213 -645 225 -611
rect 33 -651 225 -645
rect 291 -611 483 -605
rect 291 -645 303 -611
rect 471 -645 483 -611
rect 291 -651 483 -645
rect 549 -611 741 -605
rect 549 -645 561 -611
rect 729 -645 741 -611
rect 549 -651 741 -645
rect 807 -611 999 -605
rect 807 -645 819 -611
rect 987 -645 999 -611
rect 807 -651 999 -645
rect 1065 -611 1257 -605
rect 1065 -645 1077 -611
rect 1245 -645 1257 -611
rect 1065 -651 1257 -645
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
