magic
tech sky130B
magscale 1 2
timestamp 1768736825
<< error_p >>
rect -3510 645 -3452 651
rect -3392 645 -3334 651
rect -3274 645 -3216 651
rect -3156 645 -3098 651
rect -3038 645 -2980 651
rect -2920 645 -2862 651
rect -2802 645 -2744 651
rect -2684 645 -2626 651
rect -2566 645 -2508 651
rect -2448 645 -2390 651
rect -2330 645 -2272 651
rect -2212 645 -2154 651
rect -2094 645 -2036 651
rect -1976 645 -1918 651
rect -1858 645 -1800 651
rect -1740 645 -1682 651
rect -1622 645 -1564 651
rect -1504 645 -1446 651
rect -1386 645 -1328 651
rect -1268 645 -1210 651
rect -1150 645 -1092 651
rect -1032 645 -974 651
rect -914 645 -856 651
rect -796 645 -738 651
rect -678 645 -620 651
rect -560 645 -502 651
rect -442 645 -384 651
rect -324 645 -266 651
rect -206 645 -148 651
rect -88 645 -30 651
rect 30 645 88 651
rect 148 645 206 651
rect 266 645 324 651
rect 384 645 442 651
rect 502 645 560 651
rect 620 645 678 651
rect 738 645 796 651
rect 856 645 914 651
rect 974 645 1032 651
rect 1092 645 1150 651
rect 1210 645 1268 651
rect 1328 645 1386 651
rect 1446 645 1504 651
rect 1564 645 1622 651
rect 1682 645 1740 651
rect 1800 645 1858 651
rect 1918 645 1976 651
rect 2036 645 2094 651
rect 2154 645 2212 651
rect 2272 645 2330 651
rect 2390 645 2448 651
rect 2508 645 2566 651
rect 2626 645 2684 651
rect 2744 645 2802 651
rect 2862 645 2920 651
rect 2980 645 3038 651
rect 3098 645 3156 651
rect 3216 645 3274 651
rect 3334 645 3392 651
rect 3452 645 3510 651
rect -3510 611 -3498 645
rect -3392 611 -3380 645
rect -3274 611 -3262 645
rect -3156 611 -3144 645
rect -3038 611 -3026 645
rect -2920 611 -2908 645
rect -2802 611 -2790 645
rect -2684 611 -2672 645
rect -2566 611 -2554 645
rect -2448 611 -2436 645
rect -2330 611 -2318 645
rect -2212 611 -2200 645
rect -2094 611 -2082 645
rect -1976 611 -1964 645
rect -1858 611 -1846 645
rect -1740 611 -1728 645
rect -1622 611 -1610 645
rect -1504 611 -1492 645
rect -1386 611 -1374 645
rect -1268 611 -1256 645
rect -1150 611 -1138 645
rect -1032 611 -1020 645
rect -914 611 -902 645
rect -796 611 -784 645
rect -678 611 -666 645
rect -560 611 -548 645
rect -442 611 -430 645
rect -324 611 -312 645
rect -206 611 -194 645
rect -88 611 -76 645
rect 30 611 42 645
rect 148 611 160 645
rect 266 611 278 645
rect 384 611 396 645
rect 502 611 514 645
rect 620 611 632 645
rect 738 611 750 645
rect 856 611 868 645
rect 974 611 986 645
rect 1092 611 1104 645
rect 1210 611 1222 645
rect 1328 611 1340 645
rect 1446 611 1458 645
rect 1564 611 1576 645
rect 1682 611 1694 645
rect 1800 611 1812 645
rect 1918 611 1930 645
rect 2036 611 2048 645
rect 2154 611 2166 645
rect 2272 611 2284 645
rect 2390 611 2402 645
rect 2508 611 2520 645
rect 2626 611 2638 645
rect 2744 611 2756 645
rect 2862 611 2874 645
rect 2980 611 2992 645
rect 3098 611 3110 645
rect 3216 611 3228 645
rect 3334 611 3346 645
rect 3452 611 3464 645
rect -3510 605 -3452 611
rect -3392 605 -3334 611
rect -3274 605 -3216 611
rect -3156 605 -3098 611
rect -3038 605 -2980 611
rect -2920 605 -2862 611
rect -2802 605 -2744 611
rect -2684 605 -2626 611
rect -2566 605 -2508 611
rect -2448 605 -2390 611
rect -2330 605 -2272 611
rect -2212 605 -2154 611
rect -2094 605 -2036 611
rect -1976 605 -1918 611
rect -1858 605 -1800 611
rect -1740 605 -1682 611
rect -1622 605 -1564 611
rect -1504 605 -1446 611
rect -1386 605 -1328 611
rect -1268 605 -1210 611
rect -1150 605 -1092 611
rect -1032 605 -974 611
rect -914 605 -856 611
rect -796 605 -738 611
rect -678 605 -620 611
rect -560 605 -502 611
rect -442 605 -384 611
rect -324 605 -266 611
rect -206 605 -148 611
rect -88 605 -30 611
rect 30 605 88 611
rect 148 605 206 611
rect 266 605 324 611
rect 384 605 442 611
rect 502 605 560 611
rect 620 605 678 611
rect 738 605 796 611
rect 856 605 914 611
rect 974 605 1032 611
rect 1092 605 1150 611
rect 1210 605 1268 611
rect 1328 605 1386 611
rect 1446 605 1504 611
rect 1564 605 1622 611
rect 1682 605 1740 611
rect 1800 605 1858 611
rect 1918 605 1976 611
rect 2036 605 2094 611
rect 2154 605 2212 611
rect 2272 605 2330 611
rect 2390 605 2448 611
rect 2508 605 2566 611
rect 2626 605 2684 611
rect 2744 605 2802 611
rect 2862 605 2920 611
rect 2980 605 3038 611
rect 3098 605 3156 611
rect 3216 605 3274 611
rect 3334 605 3392 611
rect 3452 605 3510 611
<< nwell >>
rect -3605 -698 3605 664
<< pmos >>
rect -3511 -636 -3451 564
rect -3393 -636 -3333 564
rect -3275 -636 -3215 564
rect -3157 -636 -3097 564
rect -3039 -636 -2979 564
rect -2921 -636 -2861 564
rect -2803 -636 -2743 564
rect -2685 -636 -2625 564
rect -2567 -636 -2507 564
rect -2449 -636 -2389 564
rect -2331 -636 -2271 564
rect -2213 -636 -2153 564
rect -2095 -636 -2035 564
rect -1977 -636 -1917 564
rect -1859 -636 -1799 564
rect -1741 -636 -1681 564
rect -1623 -636 -1563 564
rect -1505 -636 -1445 564
rect -1387 -636 -1327 564
rect -1269 -636 -1209 564
rect -1151 -636 -1091 564
rect -1033 -636 -973 564
rect -915 -636 -855 564
rect -797 -636 -737 564
rect -679 -636 -619 564
rect -561 -636 -501 564
rect -443 -636 -383 564
rect -325 -636 -265 564
rect -207 -636 -147 564
rect -89 -636 -29 564
rect 29 -636 89 564
rect 147 -636 207 564
rect 265 -636 325 564
rect 383 -636 443 564
rect 501 -636 561 564
rect 619 -636 679 564
rect 737 -636 797 564
rect 855 -636 915 564
rect 973 -636 1033 564
rect 1091 -636 1151 564
rect 1209 -636 1269 564
rect 1327 -636 1387 564
rect 1445 -636 1505 564
rect 1563 -636 1623 564
rect 1681 -636 1741 564
rect 1799 -636 1859 564
rect 1917 -636 1977 564
rect 2035 -636 2095 564
rect 2153 -636 2213 564
rect 2271 -636 2331 564
rect 2389 -636 2449 564
rect 2507 -636 2567 564
rect 2625 -636 2685 564
rect 2743 -636 2803 564
rect 2861 -636 2921 564
rect 2979 -636 3039 564
rect 3097 -636 3157 564
rect 3215 -636 3275 564
rect 3333 -636 3393 564
rect 3451 -636 3511 564
<< pdiff >>
rect -3569 552 -3511 564
rect -3569 -624 -3557 552
rect -3523 -624 -3511 552
rect -3569 -636 -3511 -624
rect -3451 552 -3393 564
rect -3451 -624 -3439 552
rect -3405 -624 -3393 552
rect -3451 -636 -3393 -624
rect -3333 552 -3275 564
rect -3333 -624 -3321 552
rect -3287 -624 -3275 552
rect -3333 -636 -3275 -624
rect -3215 552 -3157 564
rect -3215 -624 -3203 552
rect -3169 -624 -3157 552
rect -3215 -636 -3157 -624
rect -3097 552 -3039 564
rect -3097 -624 -3085 552
rect -3051 -624 -3039 552
rect -3097 -636 -3039 -624
rect -2979 552 -2921 564
rect -2979 -624 -2967 552
rect -2933 -624 -2921 552
rect -2979 -636 -2921 -624
rect -2861 552 -2803 564
rect -2861 -624 -2849 552
rect -2815 -624 -2803 552
rect -2861 -636 -2803 -624
rect -2743 552 -2685 564
rect -2743 -624 -2731 552
rect -2697 -624 -2685 552
rect -2743 -636 -2685 -624
rect -2625 552 -2567 564
rect -2625 -624 -2613 552
rect -2579 -624 -2567 552
rect -2625 -636 -2567 -624
rect -2507 552 -2449 564
rect -2507 -624 -2495 552
rect -2461 -624 -2449 552
rect -2507 -636 -2449 -624
rect -2389 552 -2331 564
rect -2389 -624 -2377 552
rect -2343 -624 -2331 552
rect -2389 -636 -2331 -624
rect -2271 552 -2213 564
rect -2271 -624 -2259 552
rect -2225 -624 -2213 552
rect -2271 -636 -2213 -624
rect -2153 552 -2095 564
rect -2153 -624 -2141 552
rect -2107 -624 -2095 552
rect -2153 -636 -2095 -624
rect -2035 552 -1977 564
rect -2035 -624 -2023 552
rect -1989 -624 -1977 552
rect -2035 -636 -1977 -624
rect -1917 552 -1859 564
rect -1917 -624 -1905 552
rect -1871 -624 -1859 552
rect -1917 -636 -1859 -624
rect -1799 552 -1741 564
rect -1799 -624 -1787 552
rect -1753 -624 -1741 552
rect -1799 -636 -1741 -624
rect -1681 552 -1623 564
rect -1681 -624 -1669 552
rect -1635 -624 -1623 552
rect -1681 -636 -1623 -624
rect -1563 552 -1505 564
rect -1563 -624 -1551 552
rect -1517 -624 -1505 552
rect -1563 -636 -1505 -624
rect -1445 552 -1387 564
rect -1445 -624 -1433 552
rect -1399 -624 -1387 552
rect -1445 -636 -1387 -624
rect -1327 552 -1269 564
rect -1327 -624 -1315 552
rect -1281 -624 -1269 552
rect -1327 -636 -1269 -624
rect -1209 552 -1151 564
rect -1209 -624 -1197 552
rect -1163 -624 -1151 552
rect -1209 -636 -1151 -624
rect -1091 552 -1033 564
rect -1091 -624 -1079 552
rect -1045 -624 -1033 552
rect -1091 -636 -1033 -624
rect -973 552 -915 564
rect -973 -624 -961 552
rect -927 -624 -915 552
rect -973 -636 -915 -624
rect -855 552 -797 564
rect -855 -624 -843 552
rect -809 -624 -797 552
rect -855 -636 -797 -624
rect -737 552 -679 564
rect -737 -624 -725 552
rect -691 -624 -679 552
rect -737 -636 -679 -624
rect -619 552 -561 564
rect -619 -624 -607 552
rect -573 -624 -561 552
rect -619 -636 -561 -624
rect -501 552 -443 564
rect -501 -624 -489 552
rect -455 -624 -443 552
rect -501 -636 -443 -624
rect -383 552 -325 564
rect -383 -624 -371 552
rect -337 -624 -325 552
rect -383 -636 -325 -624
rect -265 552 -207 564
rect -265 -624 -253 552
rect -219 -624 -207 552
rect -265 -636 -207 -624
rect -147 552 -89 564
rect -147 -624 -135 552
rect -101 -624 -89 552
rect -147 -636 -89 -624
rect -29 552 29 564
rect -29 -624 -17 552
rect 17 -624 29 552
rect -29 -636 29 -624
rect 89 552 147 564
rect 89 -624 101 552
rect 135 -624 147 552
rect 89 -636 147 -624
rect 207 552 265 564
rect 207 -624 219 552
rect 253 -624 265 552
rect 207 -636 265 -624
rect 325 552 383 564
rect 325 -624 337 552
rect 371 -624 383 552
rect 325 -636 383 -624
rect 443 552 501 564
rect 443 -624 455 552
rect 489 -624 501 552
rect 443 -636 501 -624
rect 561 552 619 564
rect 561 -624 573 552
rect 607 -624 619 552
rect 561 -636 619 -624
rect 679 552 737 564
rect 679 -624 691 552
rect 725 -624 737 552
rect 679 -636 737 -624
rect 797 552 855 564
rect 797 -624 809 552
rect 843 -624 855 552
rect 797 -636 855 -624
rect 915 552 973 564
rect 915 -624 927 552
rect 961 -624 973 552
rect 915 -636 973 -624
rect 1033 552 1091 564
rect 1033 -624 1045 552
rect 1079 -624 1091 552
rect 1033 -636 1091 -624
rect 1151 552 1209 564
rect 1151 -624 1163 552
rect 1197 -624 1209 552
rect 1151 -636 1209 -624
rect 1269 552 1327 564
rect 1269 -624 1281 552
rect 1315 -624 1327 552
rect 1269 -636 1327 -624
rect 1387 552 1445 564
rect 1387 -624 1399 552
rect 1433 -624 1445 552
rect 1387 -636 1445 -624
rect 1505 552 1563 564
rect 1505 -624 1517 552
rect 1551 -624 1563 552
rect 1505 -636 1563 -624
rect 1623 552 1681 564
rect 1623 -624 1635 552
rect 1669 -624 1681 552
rect 1623 -636 1681 -624
rect 1741 552 1799 564
rect 1741 -624 1753 552
rect 1787 -624 1799 552
rect 1741 -636 1799 -624
rect 1859 552 1917 564
rect 1859 -624 1871 552
rect 1905 -624 1917 552
rect 1859 -636 1917 -624
rect 1977 552 2035 564
rect 1977 -624 1989 552
rect 2023 -624 2035 552
rect 1977 -636 2035 -624
rect 2095 552 2153 564
rect 2095 -624 2107 552
rect 2141 -624 2153 552
rect 2095 -636 2153 -624
rect 2213 552 2271 564
rect 2213 -624 2225 552
rect 2259 -624 2271 552
rect 2213 -636 2271 -624
rect 2331 552 2389 564
rect 2331 -624 2343 552
rect 2377 -624 2389 552
rect 2331 -636 2389 -624
rect 2449 552 2507 564
rect 2449 -624 2461 552
rect 2495 -624 2507 552
rect 2449 -636 2507 -624
rect 2567 552 2625 564
rect 2567 -624 2579 552
rect 2613 -624 2625 552
rect 2567 -636 2625 -624
rect 2685 552 2743 564
rect 2685 -624 2697 552
rect 2731 -624 2743 552
rect 2685 -636 2743 -624
rect 2803 552 2861 564
rect 2803 -624 2815 552
rect 2849 -624 2861 552
rect 2803 -636 2861 -624
rect 2921 552 2979 564
rect 2921 -624 2933 552
rect 2967 -624 2979 552
rect 2921 -636 2979 -624
rect 3039 552 3097 564
rect 3039 -624 3051 552
rect 3085 -624 3097 552
rect 3039 -636 3097 -624
rect 3157 552 3215 564
rect 3157 -624 3169 552
rect 3203 -624 3215 552
rect 3157 -636 3215 -624
rect 3275 552 3333 564
rect 3275 -624 3287 552
rect 3321 -624 3333 552
rect 3275 -636 3333 -624
rect 3393 552 3451 564
rect 3393 -624 3405 552
rect 3439 -624 3451 552
rect 3393 -636 3451 -624
rect 3511 552 3569 564
rect 3511 -624 3523 552
rect 3557 -624 3569 552
rect 3511 -636 3569 -624
<< pdiffc >>
rect -3557 -624 -3523 552
rect -3439 -624 -3405 552
rect -3321 -624 -3287 552
rect -3203 -624 -3169 552
rect -3085 -624 -3051 552
rect -2967 -624 -2933 552
rect -2849 -624 -2815 552
rect -2731 -624 -2697 552
rect -2613 -624 -2579 552
rect -2495 -624 -2461 552
rect -2377 -624 -2343 552
rect -2259 -624 -2225 552
rect -2141 -624 -2107 552
rect -2023 -624 -1989 552
rect -1905 -624 -1871 552
rect -1787 -624 -1753 552
rect -1669 -624 -1635 552
rect -1551 -624 -1517 552
rect -1433 -624 -1399 552
rect -1315 -624 -1281 552
rect -1197 -624 -1163 552
rect -1079 -624 -1045 552
rect -961 -624 -927 552
rect -843 -624 -809 552
rect -725 -624 -691 552
rect -607 -624 -573 552
rect -489 -624 -455 552
rect -371 -624 -337 552
rect -253 -624 -219 552
rect -135 -624 -101 552
rect -17 -624 17 552
rect 101 -624 135 552
rect 219 -624 253 552
rect 337 -624 371 552
rect 455 -624 489 552
rect 573 -624 607 552
rect 691 -624 725 552
rect 809 -624 843 552
rect 927 -624 961 552
rect 1045 -624 1079 552
rect 1163 -624 1197 552
rect 1281 -624 1315 552
rect 1399 -624 1433 552
rect 1517 -624 1551 552
rect 1635 -624 1669 552
rect 1753 -624 1787 552
rect 1871 -624 1905 552
rect 1989 -624 2023 552
rect 2107 -624 2141 552
rect 2225 -624 2259 552
rect 2343 -624 2377 552
rect 2461 -624 2495 552
rect 2579 -624 2613 552
rect 2697 -624 2731 552
rect 2815 -624 2849 552
rect 2933 -624 2967 552
rect 3051 -624 3085 552
rect 3169 -624 3203 552
rect 3287 -624 3321 552
rect 3405 -624 3439 552
rect 3523 -624 3557 552
<< poly >>
rect -3514 645 -3448 661
rect -3514 611 -3498 645
rect -3464 611 -3448 645
rect -3514 595 -3448 611
rect -3396 645 -3330 661
rect -3396 611 -3380 645
rect -3346 611 -3330 645
rect -3396 595 -3330 611
rect -3278 645 -3212 661
rect -3278 611 -3262 645
rect -3228 611 -3212 645
rect -3278 595 -3212 611
rect -3160 645 -3094 661
rect -3160 611 -3144 645
rect -3110 611 -3094 645
rect -3160 595 -3094 611
rect -3042 645 -2976 661
rect -3042 611 -3026 645
rect -2992 611 -2976 645
rect -3042 595 -2976 611
rect -2924 645 -2858 661
rect -2924 611 -2908 645
rect -2874 611 -2858 645
rect -2924 595 -2858 611
rect -2806 645 -2740 661
rect -2806 611 -2790 645
rect -2756 611 -2740 645
rect -2806 595 -2740 611
rect -2688 645 -2622 661
rect -2688 611 -2672 645
rect -2638 611 -2622 645
rect -2688 595 -2622 611
rect -2570 645 -2504 661
rect -2570 611 -2554 645
rect -2520 611 -2504 645
rect -2570 595 -2504 611
rect -2452 645 -2386 661
rect -2452 611 -2436 645
rect -2402 611 -2386 645
rect -2452 595 -2386 611
rect -2334 645 -2268 661
rect -2334 611 -2318 645
rect -2284 611 -2268 645
rect -2334 595 -2268 611
rect -2216 645 -2150 661
rect -2216 611 -2200 645
rect -2166 611 -2150 645
rect -2216 595 -2150 611
rect -2098 645 -2032 661
rect -2098 611 -2082 645
rect -2048 611 -2032 645
rect -2098 595 -2032 611
rect -1980 645 -1914 661
rect -1980 611 -1964 645
rect -1930 611 -1914 645
rect -1980 595 -1914 611
rect -1862 645 -1796 661
rect -1862 611 -1846 645
rect -1812 611 -1796 645
rect -1862 595 -1796 611
rect -1744 645 -1678 661
rect -1744 611 -1728 645
rect -1694 611 -1678 645
rect -1744 595 -1678 611
rect -1626 645 -1560 661
rect -1626 611 -1610 645
rect -1576 611 -1560 645
rect -1626 595 -1560 611
rect -1508 645 -1442 661
rect -1508 611 -1492 645
rect -1458 611 -1442 645
rect -1508 595 -1442 611
rect -1390 645 -1324 661
rect -1390 611 -1374 645
rect -1340 611 -1324 645
rect -1390 595 -1324 611
rect -1272 645 -1206 661
rect -1272 611 -1256 645
rect -1222 611 -1206 645
rect -1272 595 -1206 611
rect -1154 645 -1088 661
rect -1154 611 -1138 645
rect -1104 611 -1088 645
rect -1154 595 -1088 611
rect -1036 645 -970 661
rect -1036 611 -1020 645
rect -986 611 -970 645
rect -1036 595 -970 611
rect -918 645 -852 661
rect -918 611 -902 645
rect -868 611 -852 645
rect -918 595 -852 611
rect -800 645 -734 661
rect -800 611 -784 645
rect -750 611 -734 645
rect -800 595 -734 611
rect -682 645 -616 661
rect -682 611 -666 645
rect -632 611 -616 645
rect -682 595 -616 611
rect -564 645 -498 661
rect -564 611 -548 645
rect -514 611 -498 645
rect -564 595 -498 611
rect -446 645 -380 661
rect -446 611 -430 645
rect -396 611 -380 645
rect -446 595 -380 611
rect -328 645 -262 661
rect -328 611 -312 645
rect -278 611 -262 645
rect -328 595 -262 611
rect -210 645 -144 661
rect -210 611 -194 645
rect -160 611 -144 645
rect -210 595 -144 611
rect -92 645 -26 661
rect -92 611 -76 645
rect -42 611 -26 645
rect -92 595 -26 611
rect 26 645 92 661
rect 26 611 42 645
rect 76 611 92 645
rect 26 595 92 611
rect 144 645 210 661
rect 144 611 160 645
rect 194 611 210 645
rect 144 595 210 611
rect 262 645 328 661
rect 262 611 278 645
rect 312 611 328 645
rect 262 595 328 611
rect 380 645 446 661
rect 380 611 396 645
rect 430 611 446 645
rect 380 595 446 611
rect 498 645 564 661
rect 498 611 514 645
rect 548 611 564 645
rect 498 595 564 611
rect 616 645 682 661
rect 616 611 632 645
rect 666 611 682 645
rect 616 595 682 611
rect 734 645 800 661
rect 734 611 750 645
rect 784 611 800 645
rect 734 595 800 611
rect 852 645 918 661
rect 852 611 868 645
rect 902 611 918 645
rect 852 595 918 611
rect 970 645 1036 661
rect 970 611 986 645
rect 1020 611 1036 645
rect 970 595 1036 611
rect 1088 645 1154 661
rect 1088 611 1104 645
rect 1138 611 1154 645
rect 1088 595 1154 611
rect 1206 645 1272 661
rect 1206 611 1222 645
rect 1256 611 1272 645
rect 1206 595 1272 611
rect 1324 645 1390 661
rect 1324 611 1340 645
rect 1374 611 1390 645
rect 1324 595 1390 611
rect 1442 645 1508 661
rect 1442 611 1458 645
rect 1492 611 1508 645
rect 1442 595 1508 611
rect 1560 645 1626 661
rect 1560 611 1576 645
rect 1610 611 1626 645
rect 1560 595 1626 611
rect 1678 645 1744 661
rect 1678 611 1694 645
rect 1728 611 1744 645
rect 1678 595 1744 611
rect 1796 645 1862 661
rect 1796 611 1812 645
rect 1846 611 1862 645
rect 1796 595 1862 611
rect 1914 645 1980 661
rect 1914 611 1930 645
rect 1964 611 1980 645
rect 1914 595 1980 611
rect 2032 645 2098 661
rect 2032 611 2048 645
rect 2082 611 2098 645
rect 2032 595 2098 611
rect 2150 645 2216 661
rect 2150 611 2166 645
rect 2200 611 2216 645
rect 2150 595 2216 611
rect 2268 645 2334 661
rect 2268 611 2284 645
rect 2318 611 2334 645
rect 2268 595 2334 611
rect 2386 645 2452 661
rect 2386 611 2402 645
rect 2436 611 2452 645
rect 2386 595 2452 611
rect 2504 645 2570 661
rect 2504 611 2520 645
rect 2554 611 2570 645
rect 2504 595 2570 611
rect 2622 645 2688 661
rect 2622 611 2638 645
rect 2672 611 2688 645
rect 2622 595 2688 611
rect 2740 645 2806 661
rect 2740 611 2756 645
rect 2790 611 2806 645
rect 2740 595 2806 611
rect 2858 645 2924 661
rect 2858 611 2874 645
rect 2908 611 2924 645
rect 2858 595 2924 611
rect 2976 645 3042 661
rect 2976 611 2992 645
rect 3026 611 3042 645
rect 2976 595 3042 611
rect 3094 645 3160 661
rect 3094 611 3110 645
rect 3144 611 3160 645
rect 3094 595 3160 611
rect 3212 645 3278 661
rect 3212 611 3228 645
rect 3262 611 3278 645
rect 3212 595 3278 611
rect 3330 645 3396 661
rect 3330 611 3346 645
rect 3380 611 3396 645
rect 3330 595 3396 611
rect 3448 645 3514 661
rect 3448 611 3464 645
rect 3498 611 3514 645
rect 3448 595 3514 611
rect -3511 564 -3451 595
rect -3393 564 -3333 595
rect -3275 564 -3215 595
rect -3157 564 -3097 595
rect -3039 564 -2979 595
rect -2921 564 -2861 595
rect -2803 564 -2743 595
rect -2685 564 -2625 595
rect -2567 564 -2507 595
rect -2449 564 -2389 595
rect -2331 564 -2271 595
rect -2213 564 -2153 595
rect -2095 564 -2035 595
rect -1977 564 -1917 595
rect -1859 564 -1799 595
rect -1741 564 -1681 595
rect -1623 564 -1563 595
rect -1505 564 -1445 595
rect -1387 564 -1327 595
rect -1269 564 -1209 595
rect -1151 564 -1091 595
rect -1033 564 -973 595
rect -915 564 -855 595
rect -797 564 -737 595
rect -679 564 -619 595
rect -561 564 -501 595
rect -443 564 -383 595
rect -325 564 -265 595
rect -207 564 -147 595
rect -89 564 -29 595
rect 29 564 89 595
rect 147 564 207 595
rect 265 564 325 595
rect 383 564 443 595
rect 501 564 561 595
rect 619 564 679 595
rect 737 564 797 595
rect 855 564 915 595
rect 973 564 1033 595
rect 1091 564 1151 595
rect 1209 564 1269 595
rect 1327 564 1387 595
rect 1445 564 1505 595
rect 1563 564 1623 595
rect 1681 564 1741 595
rect 1799 564 1859 595
rect 1917 564 1977 595
rect 2035 564 2095 595
rect 2153 564 2213 595
rect 2271 564 2331 595
rect 2389 564 2449 595
rect 2507 564 2567 595
rect 2625 564 2685 595
rect 2743 564 2803 595
rect 2861 564 2921 595
rect 2979 564 3039 595
rect 3097 564 3157 595
rect 3215 564 3275 595
rect 3333 564 3393 595
rect 3451 564 3511 595
rect -3511 -662 -3451 -636
rect -3393 -662 -3333 -636
rect -3275 -662 -3215 -636
rect -3157 -662 -3097 -636
rect -3039 -662 -2979 -636
rect -2921 -662 -2861 -636
rect -2803 -662 -2743 -636
rect -2685 -662 -2625 -636
rect -2567 -662 -2507 -636
rect -2449 -662 -2389 -636
rect -2331 -662 -2271 -636
rect -2213 -662 -2153 -636
rect -2095 -662 -2035 -636
rect -1977 -662 -1917 -636
rect -1859 -662 -1799 -636
rect -1741 -662 -1681 -636
rect -1623 -662 -1563 -636
rect -1505 -662 -1445 -636
rect -1387 -662 -1327 -636
rect -1269 -662 -1209 -636
rect -1151 -662 -1091 -636
rect -1033 -662 -973 -636
rect -915 -662 -855 -636
rect -797 -662 -737 -636
rect -679 -662 -619 -636
rect -561 -662 -501 -636
rect -443 -662 -383 -636
rect -325 -662 -265 -636
rect -207 -662 -147 -636
rect -89 -662 -29 -636
rect 29 -662 89 -636
rect 147 -662 207 -636
rect 265 -662 325 -636
rect 383 -662 443 -636
rect 501 -662 561 -636
rect 619 -662 679 -636
rect 737 -662 797 -636
rect 855 -662 915 -636
rect 973 -662 1033 -636
rect 1091 -662 1151 -636
rect 1209 -662 1269 -636
rect 1327 -662 1387 -636
rect 1445 -662 1505 -636
rect 1563 -662 1623 -636
rect 1681 -662 1741 -636
rect 1799 -662 1859 -636
rect 1917 -662 1977 -636
rect 2035 -662 2095 -636
rect 2153 -662 2213 -636
rect 2271 -662 2331 -636
rect 2389 -662 2449 -636
rect 2507 -662 2567 -636
rect 2625 -662 2685 -636
rect 2743 -662 2803 -636
rect 2861 -662 2921 -636
rect 2979 -662 3039 -636
rect 3097 -662 3157 -636
rect 3215 -662 3275 -636
rect 3333 -662 3393 -636
rect 3451 -662 3511 -636
<< polycont >>
rect -3498 611 -3464 645
rect -3380 611 -3346 645
rect -3262 611 -3228 645
rect -3144 611 -3110 645
rect -3026 611 -2992 645
rect -2908 611 -2874 645
rect -2790 611 -2756 645
rect -2672 611 -2638 645
rect -2554 611 -2520 645
rect -2436 611 -2402 645
rect -2318 611 -2284 645
rect -2200 611 -2166 645
rect -2082 611 -2048 645
rect -1964 611 -1930 645
rect -1846 611 -1812 645
rect -1728 611 -1694 645
rect -1610 611 -1576 645
rect -1492 611 -1458 645
rect -1374 611 -1340 645
rect -1256 611 -1222 645
rect -1138 611 -1104 645
rect -1020 611 -986 645
rect -902 611 -868 645
rect -784 611 -750 645
rect -666 611 -632 645
rect -548 611 -514 645
rect -430 611 -396 645
rect -312 611 -278 645
rect -194 611 -160 645
rect -76 611 -42 645
rect 42 611 76 645
rect 160 611 194 645
rect 278 611 312 645
rect 396 611 430 645
rect 514 611 548 645
rect 632 611 666 645
rect 750 611 784 645
rect 868 611 902 645
rect 986 611 1020 645
rect 1104 611 1138 645
rect 1222 611 1256 645
rect 1340 611 1374 645
rect 1458 611 1492 645
rect 1576 611 1610 645
rect 1694 611 1728 645
rect 1812 611 1846 645
rect 1930 611 1964 645
rect 2048 611 2082 645
rect 2166 611 2200 645
rect 2284 611 2318 645
rect 2402 611 2436 645
rect 2520 611 2554 645
rect 2638 611 2672 645
rect 2756 611 2790 645
rect 2874 611 2908 645
rect 2992 611 3026 645
rect 3110 611 3144 645
rect 3228 611 3262 645
rect 3346 611 3380 645
rect 3464 611 3498 645
<< locali >>
rect -3514 611 -3498 645
rect -3464 611 -3448 645
rect -3396 611 -3380 645
rect -3346 611 -3330 645
rect -3278 611 -3262 645
rect -3228 611 -3212 645
rect -3160 611 -3144 645
rect -3110 611 -3094 645
rect -3042 611 -3026 645
rect -2992 611 -2976 645
rect -2924 611 -2908 645
rect -2874 611 -2858 645
rect -2806 611 -2790 645
rect -2756 611 -2740 645
rect -2688 611 -2672 645
rect -2638 611 -2622 645
rect -2570 611 -2554 645
rect -2520 611 -2504 645
rect -2452 611 -2436 645
rect -2402 611 -2386 645
rect -2334 611 -2318 645
rect -2284 611 -2268 645
rect -2216 611 -2200 645
rect -2166 611 -2150 645
rect -2098 611 -2082 645
rect -2048 611 -2032 645
rect -1980 611 -1964 645
rect -1930 611 -1914 645
rect -1862 611 -1846 645
rect -1812 611 -1796 645
rect -1744 611 -1728 645
rect -1694 611 -1678 645
rect -1626 611 -1610 645
rect -1576 611 -1560 645
rect -1508 611 -1492 645
rect -1458 611 -1442 645
rect -1390 611 -1374 645
rect -1340 611 -1324 645
rect -1272 611 -1256 645
rect -1222 611 -1206 645
rect -1154 611 -1138 645
rect -1104 611 -1088 645
rect -1036 611 -1020 645
rect -986 611 -970 645
rect -918 611 -902 645
rect -868 611 -852 645
rect -800 611 -784 645
rect -750 611 -734 645
rect -682 611 -666 645
rect -632 611 -616 645
rect -564 611 -548 645
rect -514 611 -498 645
rect -446 611 -430 645
rect -396 611 -380 645
rect -328 611 -312 645
rect -278 611 -262 645
rect -210 611 -194 645
rect -160 611 -144 645
rect -92 611 -76 645
rect -42 611 -26 645
rect 26 611 42 645
rect 76 611 92 645
rect 144 611 160 645
rect 194 611 210 645
rect 262 611 278 645
rect 312 611 328 645
rect 380 611 396 645
rect 430 611 446 645
rect 498 611 514 645
rect 548 611 564 645
rect 616 611 632 645
rect 666 611 682 645
rect 734 611 750 645
rect 784 611 800 645
rect 852 611 868 645
rect 902 611 918 645
rect 970 611 986 645
rect 1020 611 1036 645
rect 1088 611 1104 645
rect 1138 611 1154 645
rect 1206 611 1222 645
rect 1256 611 1272 645
rect 1324 611 1340 645
rect 1374 611 1390 645
rect 1442 611 1458 645
rect 1492 611 1508 645
rect 1560 611 1576 645
rect 1610 611 1626 645
rect 1678 611 1694 645
rect 1728 611 1744 645
rect 1796 611 1812 645
rect 1846 611 1862 645
rect 1914 611 1930 645
rect 1964 611 1980 645
rect 2032 611 2048 645
rect 2082 611 2098 645
rect 2150 611 2166 645
rect 2200 611 2216 645
rect 2268 611 2284 645
rect 2318 611 2334 645
rect 2386 611 2402 645
rect 2436 611 2452 645
rect 2504 611 2520 645
rect 2554 611 2570 645
rect 2622 611 2638 645
rect 2672 611 2688 645
rect 2740 611 2756 645
rect 2790 611 2806 645
rect 2858 611 2874 645
rect 2908 611 2924 645
rect 2976 611 2992 645
rect 3026 611 3042 645
rect 3094 611 3110 645
rect 3144 611 3160 645
rect 3212 611 3228 645
rect 3262 611 3278 645
rect 3330 611 3346 645
rect 3380 611 3396 645
rect 3448 611 3464 645
rect 3498 611 3514 645
rect -3557 552 -3523 568
rect -3557 -640 -3523 -624
rect -3439 552 -3405 568
rect -3439 -640 -3405 -624
rect -3321 552 -3287 568
rect -3321 -640 -3287 -624
rect -3203 552 -3169 568
rect -3203 -640 -3169 -624
rect -3085 552 -3051 568
rect -3085 -640 -3051 -624
rect -2967 552 -2933 568
rect -2967 -640 -2933 -624
rect -2849 552 -2815 568
rect -2849 -640 -2815 -624
rect -2731 552 -2697 568
rect -2731 -640 -2697 -624
rect -2613 552 -2579 568
rect -2613 -640 -2579 -624
rect -2495 552 -2461 568
rect -2495 -640 -2461 -624
rect -2377 552 -2343 568
rect -2377 -640 -2343 -624
rect -2259 552 -2225 568
rect -2259 -640 -2225 -624
rect -2141 552 -2107 568
rect -2141 -640 -2107 -624
rect -2023 552 -1989 568
rect -2023 -640 -1989 -624
rect -1905 552 -1871 568
rect -1905 -640 -1871 -624
rect -1787 552 -1753 568
rect -1787 -640 -1753 -624
rect -1669 552 -1635 568
rect -1669 -640 -1635 -624
rect -1551 552 -1517 568
rect -1551 -640 -1517 -624
rect -1433 552 -1399 568
rect -1433 -640 -1399 -624
rect -1315 552 -1281 568
rect -1315 -640 -1281 -624
rect -1197 552 -1163 568
rect -1197 -640 -1163 -624
rect -1079 552 -1045 568
rect -1079 -640 -1045 -624
rect -961 552 -927 568
rect -961 -640 -927 -624
rect -843 552 -809 568
rect -843 -640 -809 -624
rect -725 552 -691 568
rect -725 -640 -691 -624
rect -607 552 -573 568
rect -607 -640 -573 -624
rect -489 552 -455 568
rect -489 -640 -455 -624
rect -371 552 -337 568
rect -371 -640 -337 -624
rect -253 552 -219 568
rect -253 -640 -219 -624
rect -135 552 -101 568
rect -135 -640 -101 -624
rect -17 552 17 568
rect -17 -640 17 -624
rect 101 552 135 568
rect 101 -640 135 -624
rect 219 552 253 568
rect 219 -640 253 -624
rect 337 552 371 568
rect 337 -640 371 -624
rect 455 552 489 568
rect 455 -640 489 -624
rect 573 552 607 568
rect 573 -640 607 -624
rect 691 552 725 568
rect 691 -640 725 -624
rect 809 552 843 568
rect 809 -640 843 -624
rect 927 552 961 568
rect 927 -640 961 -624
rect 1045 552 1079 568
rect 1045 -640 1079 -624
rect 1163 552 1197 568
rect 1163 -640 1197 -624
rect 1281 552 1315 568
rect 1281 -640 1315 -624
rect 1399 552 1433 568
rect 1399 -640 1433 -624
rect 1517 552 1551 568
rect 1517 -640 1551 -624
rect 1635 552 1669 568
rect 1635 -640 1669 -624
rect 1753 552 1787 568
rect 1753 -640 1787 -624
rect 1871 552 1905 568
rect 1871 -640 1905 -624
rect 1989 552 2023 568
rect 1989 -640 2023 -624
rect 2107 552 2141 568
rect 2107 -640 2141 -624
rect 2225 552 2259 568
rect 2225 -640 2259 -624
rect 2343 552 2377 568
rect 2343 -640 2377 -624
rect 2461 552 2495 568
rect 2461 -640 2495 -624
rect 2579 552 2613 568
rect 2579 -640 2613 -624
rect 2697 552 2731 568
rect 2697 -640 2731 -624
rect 2815 552 2849 568
rect 2815 -640 2849 -624
rect 2933 552 2967 568
rect 2933 -640 2967 -624
rect 3051 552 3085 568
rect 3051 -640 3085 -624
rect 3169 552 3203 568
rect 3169 -640 3203 -624
rect 3287 552 3321 568
rect 3287 -640 3321 -624
rect 3405 552 3439 568
rect 3405 -640 3439 -624
rect 3523 552 3557 568
rect 3523 -640 3557 -624
<< viali >>
rect -3498 611 -3464 645
rect -3380 611 -3346 645
rect -3262 611 -3228 645
rect -3144 611 -3110 645
rect -3026 611 -2992 645
rect -2908 611 -2874 645
rect -2790 611 -2756 645
rect -2672 611 -2638 645
rect -2554 611 -2520 645
rect -2436 611 -2402 645
rect -2318 611 -2284 645
rect -2200 611 -2166 645
rect -2082 611 -2048 645
rect -1964 611 -1930 645
rect -1846 611 -1812 645
rect -1728 611 -1694 645
rect -1610 611 -1576 645
rect -1492 611 -1458 645
rect -1374 611 -1340 645
rect -1256 611 -1222 645
rect -1138 611 -1104 645
rect -1020 611 -986 645
rect -902 611 -868 645
rect -784 611 -750 645
rect -666 611 -632 645
rect -548 611 -514 645
rect -430 611 -396 645
rect -312 611 -278 645
rect -194 611 -160 645
rect -76 611 -42 645
rect 42 611 76 645
rect 160 611 194 645
rect 278 611 312 645
rect 396 611 430 645
rect 514 611 548 645
rect 632 611 666 645
rect 750 611 784 645
rect 868 611 902 645
rect 986 611 1020 645
rect 1104 611 1138 645
rect 1222 611 1256 645
rect 1340 611 1374 645
rect 1458 611 1492 645
rect 1576 611 1610 645
rect 1694 611 1728 645
rect 1812 611 1846 645
rect 1930 611 1964 645
rect 2048 611 2082 645
rect 2166 611 2200 645
rect 2284 611 2318 645
rect 2402 611 2436 645
rect 2520 611 2554 645
rect 2638 611 2672 645
rect 2756 611 2790 645
rect 2874 611 2908 645
rect 2992 611 3026 645
rect 3110 611 3144 645
rect 3228 611 3262 645
rect 3346 611 3380 645
rect 3464 611 3498 645
rect -3557 -624 -3523 552
rect -3439 -624 -3405 552
rect -3321 -624 -3287 552
rect -3203 -624 -3169 552
rect -3085 -624 -3051 552
rect -2967 -624 -2933 552
rect -2849 -624 -2815 552
rect -2731 -624 -2697 552
rect -2613 -624 -2579 552
rect -2495 -624 -2461 552
rect -2377 -624 -2343 552
rect -2259 -624 -2225 552
rect -2141 -624 -2107 552
rect -2023 -624 -1989 552
rect -1905 -624 -1871 552
rect -1787 -624 -1753 552
rect -1669 -624 -1635 552
rect -1551 -624 -1517 552
rect -1433 -624 -1399 552
rect -1315 -624 -1281 552
rect -1197 -624 -1163 552
rect -1079 -624 -1045 552
rect -961 -624 -927 552
rect -843 -624 -809 552
rect -725 -624 -691 552
rect -607 -624 -573 552
rect -489 -624 -455 552
rect -371 -624 -337 552
rect -253 -624 -219 552
rect -135 -624 -101 552
rect -17 -624 17 552
rect 101 -624 135 552
rect 219 -624 253 552
rect 337 -624 371 552
rect 455 -624 489 552
rect 573 -624 607 552
rect 691 -624 725 552
rect 809 -624 843 552
rect 927 -624 961 552
rect 1045 -624 1079 552
rect 1163 -624 1197 552
rect 1281 -624 1315 552
rect 1399 -624 1433 552
rect 1517 -624 1551 552
rect 1635 -624 1669 552
rect 1753 -624 1787 552
rect 1871 -624 1905 552
rect 1989 -624 2023 552
rect 2107 -624 2141 552
rect 2225 -624 2259 552
rect 2343 -624 2377 552
rect 2461 -624 2495 552
rect 2579 -624 2613 552
rect 2697 -624 2731 552
rect 2815 -624 2849 552
rect 2933 -624 2967 552
rect 3051 -624 3085 552
rect 3169 -624 3203 552
rect 3287 -624 3321 552
rect 3405 -624 3439 552
rect 3523 -624 3557 552
<< metal1 >>
rect -3510 645 -3452 651
rect -3510 611 -3498 645
rect -3464 611 -3452 645
rect -3510 605 -3452 611
rect -3392 645 -3334 651
rect -3392 611 -3380 645
rect -3346 611 -3334 645
rect -3392 605 -3334 611
rect -3274 645 -3216 651
rect -3274 611 -3262 645
rect -3228 611 -3216 645
rect -3274 605 -3216 611
rect -3156 645 -3098 651
rect -3156 611 -3144 645
rect -3110 611 -3098 645
rect -3156 605 -3098 611
rect -3038 645 -2980 651
rect -3038 611 -3026 645
rect -2992 611 -2980 645
rect -3038 605 -2980 611
rect -2920 645 -2862 651
rect -2920 611 -2908 645
rect -2874 611 -2862 645
rect -2920 605 -2862 611
rect -2802 645 -2744 651
rect -2802 611 -2790 645
rect -2756 611 -2744 645
rect -2802 605 -2744 611
rect -2684 645 -2626 651
rect -2684 611 -2672 645
rect -2638 611 -2626 645
rect -2684 605 -2626 611
rect -2566 645 -2508 651
rect -2566 611 -2554 645
rect -2520 611 -2508 645
rect -2566 605 -2508 611
rect -2448 645 -2390 651
rect -2448 611 -2436 645
rect -2402 611 -2390 645
rect -2448 605 -2390 611
rect -2330 645 -2272 651
rect -2330 611 -2318 645
rect -2284 611 -2272 645
rect -2330 605 -2272 611
rect -2212 645 -2154 651
rect -2212 611 -2200 645
rect -2166 611 -2154 645
rect -2212 605 -2154 611
rect -2094 645 -2036 651
rect -2094 611 -2082 645
rect -2048 611 -2036 645
rect -2094 605 -2036 611
rect -1976 645 -1918 651
rect -1976 611 -1964 645
rect -1930 611 -1918 645
rect -1976 605 -1918 611
rect -1858 645 -1800 651
rect -1858 611 -1846 645
rect -1812 611 -1800 645
rect -1858 605 -1800 611
rect -1740 645 -1682 651
rect -1740 611 -1728 645
rect -1694 611 -1682 645
rect -1740 605 -1682 611
rect -1622 645 -1564 651
rect -1622 611 -1610 645
rect -1576 611 -1564 645
rect -1622 605 -1564 611
rect -1504 645 -1446 651
rect -1504 611 -1492 645
rect -1458 611 -1446 645
rect -1504 605 -1446 611
rect -1386 645 -1328 651
rect -1386 611 -1374 645
rect -1340 611 -1328 645
rect -1386 605 -1328 611
rect -1268 645 -1210 651
rect -1268 611 -1256 645
rect -1222 611 -1210 645
rect -1268 605 -1210 611
rect -1150 645 -1092 651
rect -1150 611 -1138 645
rect -1104 611 -1092 645
rect -1150 605 -1092 611
rect -1032 645 -974 651
rect -1032 611 -1020 645
rect -986 611 -974 645
rect -1032 605 -974 611
rect -914 645 -856 651
rect -914 611 -902 645
rect -868 611 -856 645
rect -914 605 -856 611
rect -796 645 -738 651
rect -796 611 -784 645
rect -750 611 -738 645
rect -796 605 -738 611
rect -678 645 -620 651
rect -678 611 -666 645
rect -632 611 -620 645
rect -678 605 -620 611
rect -560 645 -502 651
rect -560 611 -548 645
rect -514 611 -502 645
rect -560 605 -502 611
rect -442 645 -384 651
rect -442 611 -430 645
rect -396 611 -384 645
rect -442 605 -384 611
rect -324 645 -266 651
rect -324 611 -312 645
rect -278 611 -266 645
rect -324 605 -266 611
rect -206 645 -148 651
rect -206 611 -194 645
rect -160 611 -148 645
rect -206 605 -148 611
rect -88 645 -30 651
rect -88 611 -76 645
rect -42 611 -30 645
rect -88 605 -30 611
rect 30 645 88 651
rect 30 611 42 645
rect 76 611 88 645
rect 30 605 88 611
rect 148 645 206 651
rect 148 611 160 645
rect 194 611 206 645
rect 148 605 206 611
rect 266 645 324 651
rect 266 611 278 645
rect 312 611 324 645
rect 266 605 324 611
rect 384 645 442 651
rect 384 611 396 645
rect 430 611 442 645
rect 384 605 442 611
rect 502 645 560 651
rect 502 611 514 645
rect 548 611 560 645
rect 502 605 560 611
rect 620 645 678 651
rect 620 611 632 645
rect 666 611 678 645
rect 620 605 678 611
rect 738 645 796 651
rect 738 611 750 645
rect 784 611 796 645
rect 738 605 796 611
rect 856 645 914 651
rect 856 611 868 645
rect 902 611 914 645
rect 856 605 914 611
rect 974 645 1032 651
rect 974 611 986 645
rect 1020 611 1032 645
rect 974 605 1032 611
rect 1092 645 1150 651
rect 1092 611 1104 645
rect 1138 611 1150 645
rect 1092 605 1150 611
rect 1210 645 1268 651
rect 1210 611 1222 645
rect 1256 611 1268 645
rect 1210 605 1268 611
rect 1328 645 1386 651
rect 1328 611 1340 645
rect 1374 611 1386 645
rect 1328 605 1386 611
rect 1446 645 1504 651
rect 1446 611 1458 645
rect 1492 611 1504 645
rect 1446 605 1504 611
rect 1564 645 1622 651
rect 1564 611 1576 645
rect 1610 611 1622 645
rect 1564 605 1622 611
rect 1682 645 1740 651
rect 1682 611 1694 645
rect 1728 611 1740 645
rect 1682 605 1740 611
rect 1800 645 1858 651
rect 1800 611 1812 645
rect 1846 611 1858 645
rect 1800 605 1858 611
rect 1918 645 1976 651
rect 1918 611 1930 645
rect 1964 611 1976 645
rect 1918 605 1976 611
rect 2036 645 2094 651
rect 2036 611 2048 645
rect 2082 611 2094 645
rect 2036 605 2094 611
rect 2154 645 2212 651
rect 2154 611 2166 645
rect 2200 611 2212 645
rect 2154 605 2212 611
rect 2272 645 2330 651
rect 2272 611 2284 645
rect 2318 611 2330 645
rect 2272 605 2330 611
rect 2390 645 2448 651
rect 2390 611 2402 645
rect 2436 611 2448 645
rect 2390 605 2448 611
rect 2508 645 2566 651
rect 2508 611 2520 645
rect 2554 611 2566 645
rect 2508 605 2566 611
rect 2626 645 2684 651
rect 2626 611 2638 645
rect 2672 611 2684 645
rect 2626 605 2684 611
rect 2744 645 2802 651
rect 2744 611 2756 645
rect 2790 611 2802 645
rect 2744 605 2802 611
rect 2862 645 2920 651
rect 2862 611 2874 645
rect 2908 611 2920 645
rect 2862 605 2920 611
rect 2980 645 3038 651
rect 2980 611 2992 645
rect 3026 611 3038 645
rect 2980 605 3038 611
rect 3098 645 3156 651
rect 3098 611 3110 645
rect 3144 611 3156 645
rect 3098 605 3156 611
rect 3216 645 3274 651
rect 3216 611 3228 645
rect 3262 611 3274 645
rect 3216 605 3274 611
rect 3334 645 3392 651
rect 3334 611 3346 645
rect 3380 611 3392 645
rect 3334 605 3392 611
rect 3452 645 3510 651
rect 3452 611 3464 645
rect 3498 611 3510 645
rect 3452 605 3510 611
rect -3563 552 -3517 564
rect -3563 -624 -3557 552
rect -3523 -624 -3517 552
rect -3563 -636 -3517 -624
rect -3445 552 -3399 564
rect -3445 -624 -3439 552
rect -3405 -624 -3399 552
rect -3445 -636 -3399 -624
rect -3327 552 -3281 564
rect -3327 -624 -3321 552
rect -3287 -624 -3281 552
rect -3327 -636 -3281 -624
rect -3209 552 -3163 564
rect -3209 -624 -3203 552
rect -3169 -624 -3163 552
rect -3209 -636 -3163 -624
rect -3091 552 -3045 564
rect -3091 -624 -3085 552
rect -3051 -624 -3045 552
rect -3091 -636 -3045 -624
rect -2973 552 -2927 564
rect -2973 -624 -2967 552
rect -2933 -624 -2927 552
rect -2973 -636 -2927 -624
rect -2855 552 -2809 564
rect -2855 -624 -2849 552
rect -2815 -624 -2809 552
rect -2855 -636 -2809 -624
rect -2737 552 -2691 564
rect -2737 -624 -2731 552
rect -2697 -624 -2691 552
rect -2737 -636 -2691 -624
rect -2619 552 -2573 564
rect -2619 -624 -2613 552
rect -2579 -624 -2573 552
rect -2619 -636 -2573 -624
rect -2501 552 -2455 564
rect -2501 -624 -2495 552
rect -2461 -624 -2455 552
rect -2501 -636 -2455 -624
rect -2383 552 -2337 564
rect -2383 -624 -2377 552
rect -2343 -624 -2337 552
rect -2383 -636 -2337 -624
rect -2265 552 -2219 564
rect -2265 -624 -2259 552
rect -2225 -624 -2219 552
rect -2265 -636 -2219 -624
rect -2147 552 -2101 564
rect -2147 -624 -2141 552
rect -2107 -624 -2101 552
rect -2147 -636 -2101 -624
rect -2029 552 -1983 564
rect -2029 -624 -2023 552
rect -1989 -624 -1983 552
rect -2029 -636 -1983 -624
rect -1911 552 -1865 564
rect -1911 -624 -1905 552
rect -1871 -624 -1865 552
rect -1911 -636 -1865 -624
rect -1793 552 -1747 564
rect -1793 -624 -1787 552
rect -1753 -624 -1747 552
rect -1793 -636 -1747 -624
rect -1675 552 -1629 564
rect -1675 -624 -1669 552
rect -1635 -624 -1629 552
rect -1675 -636 -1629 -624
rect -1557 552 -1511 564
rect -1557 -624 -1551 552
rect -1517 -624 -1511 552
rect -1557 -636 -1511 -624
rect -1439 552 -1393 564
rect -1439 -624 -1433 552
rect -1399 -624 -1393 552
rect -1439 -636 -1393 -624
rect -1321 552 -1275 564
rect -1321 -624 -1315 552
rect -1281 -624 -1275 552
rect -1321 -636 -1275 -624
rect -1203 552 -1157 564
rect -1203 -624 -1197 552
rect -1163 -624 -1157 552
rect -1203 -636 -1157 -624
rect -1085 552 -1039 564
rect -1085 -624 -1079 552
rect -1045 -624 -1039 552
rect -1085 -636 -1039 -624
rect -967 552 -921 564
rect -967 -624 -961 552
rect -927 -624 -921 552
rect -967 -636 -921 -624
rect -849 552 -803 564
rect -849 -624 -843 552
rect -809 -624 -803 552
rect -849 -636 -803 -624
rect -731 552 -685 564
rect -731 -624 -725 552
rect -691 -624 -685 552
rect -731 -636 -685 -624
rect -613 552 -567 564
rect -613 -624 -607 552
rect -573 -624 -567 552
rect -613 -636 -567 -624
rect -495 552 -449 564
rect -495 -624 -489 552
rect -455 -624 -449 552
rect -495 -636 -449 -624
rect -377 552 -331 564
rect -377 -624 -371 552
rect -337 -624 -331 552
rect -377 -636 -331 -624
rect -259 552 -213 564
rect -259 -624 -253 552
rect -219 -624 -213 552
rect -259 -636 -213 -624
rect -141 552 -95 564
rect -141 -624 -135 552
rect -101 -624 -95 552
rect -141 -636 -95 -624
rect -23 552 23 564
rect -23 -624 -17 552
rect 17 -624 23 552
rect -23 -636 23 -624
rect 95 552 141 564
rect 95 -624 101 552
rect 135 -624 141 552
rect 95 -636 141 -624
rect 213 552 259 564
rect 213 -624 219 552
rect 253 -624 259 552
rect 213 -636 259 -624
rect 331 552 377 564
rect 331 -624 337 552
rect 371 -624 377 552
rect 331 -636 377 -624
rect 449 552 495 564
rect 449 -624 455 552
rect 489 -624 495 552
rect 449 -636 495 -624
rect 567 552 613 564
rect 567 -624 573 552
rect 607 -624 613 552
rect 567 -636 613 -624
rect 685 552 731 564
rect 685 -624 691 552
rect 725 -624 731 552
rect 685 -636 731 -624
rect 803 552 849 564
rect 803 -624 809 552
rect 843 -624 849 552
rect 803 -636 849 -624
rect 921 552 967 564
rect 921 -624 927 552
rect 961 -624 967 552
rect 921 -636 967 -624
rect 1039 552 1085 564
rect 1039 -624 1045 552
rect 1079 -624 1085 552
rect 1039 -636 1085 -624
rect 1157 552 1203 564
rect 1157 -624 1163 552
rect 1197 -624 1203 552
rect 1157 -636 1203 -624
rect 1275 552 1321 564
rect 1275 -624 1281 552
rect 1315 -624 1321 552
rect 1275 -636 1321 -624
rect 1393 552 1439 564
rect 1393 -624 1399 552
rect 1433 -624 1439 552
rect 1393 -636 1439 -624
rect 1511 552 1557 564
rect 1511 -624 1517 552
rect 1551 -624 1557 552
rect 1511 -636 1557 -624
rect 1629 552 1675 564
rect 1629 -624 1635 552
rect 1669 -624 1675 552
rect 1629 -636 1675 -624
rect 1747 552 1793 564
rect 1747 -624 1753 552
rect 1787 -624 1793 552
rect 1747 -636 1793 -624
rect 1865 552 1911 564
rect 1865 -624 1871 552
rect 1905 -624 1911 552
rect 1865 -636 1911 -624
rect 1983 552 2029 564
rect 1983 -624 1989 552
rect 2023 -624 2029 552
rect 1983 -636 2029 -624
rect 2101 552 2147 564
rect 2101 -624 2107 552
rect 2141 -624 2147 552
rect 2101 -636 2147 -624
rect 2219 552 2265 564
rect 2219 -624 2225 552
rect 2259 -624 2265 552
rect 2219 -636 2265 -624
rect 2337 552 2383 564
rect 2337 -624 2343 552
rect 2377 -624 2383 552
rect 2337 -636 2383 -624
rect 2455 552 2501 564
rect 2455 -624 2461 552
rect 2495 -624 2501 552
rect 2455 -636 2501 -624
rect 2573 552 2619 564
rect 2573 -624 2579 552
rect 2613 -624 2619 552
rect 2573 -636 2619 -624
rect 2691 552 2737 564
rect 2691 -624 2697 552
rect 2731 -624 2737 552
rect 2691 -636 2737 -624
rect 2809 552 2855 564
rect 2809 -624 2815 552
rect 2849 -624 2855 552
rect 2809 -636 2855 -624
rect 2927 552 2973 564
rect 2927 -624 2933 552
rect 2967 -624 2973 552
rect 2927 -636 2973 -624
rect 3045 552 3091 564
rect 3045 -624 3051 552
rect 3085 -624 3091 552
rect 3045 -636 3091 -624
rect 3163 552 3209 564
rect 3163 -624 3169 552
rect 3203 -624 3209 552
rect 3163 -636 3209 -624
rect 3281 552 3327 564
rect 3281 -624 3287 552
rect 3321 -624 3327 552
rect 3281 -636 3327 -624
rect 3399 552 3445 564
rect 3399 -624 3405 552
rect 3439 -624 3445 552
rect 3399 -636 3445 -624
rect 3517 552 3563 564
rect 3517 -624 3523 552
rect 3557 -624 3563 552
rect 3517 -636 3563 -624
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.3 m 1 nf 60 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
