VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mete_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_mete_opamp ;
  ORIGIN 13.100 -26.490 ;
  SIZE 46.220 BY 37.510 ;
  PIN Vin-
    ANTENNAGATEAREA 17.010000 ;
    PORT
      LAYER li1 ;
        RECT -12.520 47.170 -12.350 48.170 ;
        RECT -12.520 45.880 -12.350 46.880 ;
        RECT -12.520 44.590 -12.350 45.590 ;
      LAYER mcon ;
        RECT -12.520 47.250 -12.350 48.090 ;
        RECT -12.520 45.960 -12.350 46.800 ;
        RECT -12.520 44.670 -12.350 45.510 ;
      LAYER met1 ;
        RECT -12.830 44.590 -12.300 48.200 ;
        RECT -12.830 43.780 -12.350 44.590 ;
        RECT -12.830 43.000 -10.900 43.780 ;
    END
  END Vin-
  PIN Vin+
    ANTENNAGATEAREA 17.010000 ;
    PORT
      LAYER li1 ;
        RECT 0.990 47.170 1.160 48.170 ;
        RECT 0.990 45.880 1.160 46.880 ;
        RECT 0.990 44.590 1.160 45.590 ;
      LAYER mcon ;
        RECT 0.990 47.250 1.160 48.090 ;
        RECT 0.990 45.960 1.160 46.800 ;
        RECT 0.990 44.670 1.160 45.510 ;
      LAYER met1 ;
        RECT 0.960 47.900 1.190 48.150 ;
        RECT 0.900 47.270 1.210 47.900 ;
        RECT 0.960 46.900 1.210 47.270 ;
        RECT 0.940 46.800 2.400 46.900 ;
        RECT 0.900 46.000 2.400 46.800 ;
        RECT 0.900 45.980 1.210 46.000 ;
        RECT 0.960 45.500 1.210 45.980 ;
        RECT 0.900 44.700 1.210 45.500 ;
        RECT 0.960 44.610 1.190 44.700 ;
    END
  END Vin+
  PIN Ptatin
    ANTENNAGATEAREA 65.150002 ;
    ANTENNADIFFAREA 3.190000 ;
    PORT
      LAYER li1 ;
        RECT 19.000 60.920 19.170 61.920 ;
        RECT 19.000 59.630 19.170 60.630 ;
        RECT 19.000 58.340 19.170 59.340 ;
        RECT 11.385 56.770 11.555 57.100 ;
        RECT 19.000 57.050 19.170 58.050 ;
        RECT 11.770 56.630 12.810 56.800 ;
        RECT 19.000 55.760 19.170 56.760 ;
        RECT 3.380 53.390 3.550 54.390 ;
        RECT 8.930 53.390 9.100 54.390 ;
        RECT 11.570 54.190 11.740 55.190 ;
        RECT 11.910 53.960 16.950 54.130 ;
        RECT 11.920 53.350 16.960 53.520 ;
        RECT 11.580 52.290 11.750 53.290 ;
        RECT 0.820 42.660 0.990 43.660 ;
        RECT 0.820 41.370 0.990 42.370 ;
        RECT 0.820 40.080 0.990 41.080 ;
        RECT 0.820 38.790 0.990 39.790 ;
      LAYER mcon ;
        RECT 19.000 61.000 19.170 61.840 ;
        RECT 19.000 59.710 19.170 60.550 ;
        RECT 19.000 58.420 19.170 59.260 ;
        RECT 19.000 57.130 19.170 57.970 ;
        RECT 11.385 56.850 11.555 57.020 ;
        RECT 11.850 56.630 12.730 56.800 ;
        RECT 19.000 55.840 19.170 56.680 ;
        RECT 3.380 53.470 3.550 54.310 ;
        RECT 8.930 53.470 9.100 54.310 ;
        RECT 11.570 54.270 11.740 55.110 ;
        RECT 11.990 53.960 16.870 54.130 ;
        RECT 12.000 53.350 16.880 53.520 ;
        RECT 11.580 52.370 11.750 53.210 ;
        RECT 0.820 42.740 0.990 43.580 ;
        RECT 0.820 41.450 0.990 42.290 ;
        RECT 0.820 40.160 0.990 41.000 ;
        RECT 0.820 38.870 0.990 39.710 ;
      LAYER met1 ;
        RECT 18.850 58.400 19.200 61.900 ;
        RECT 18.100 57.400 19.200 58.400 ;
        RECT 10.900 56.640 11.600 57.100 ;
        RECT 11.790 56.800 12.790 56.830 ;
        RECT 11.740 56.640 12.810 56.800 ;
        RECT 10.900 56.400 12.810 56.640 ;
        RECT 10.900 55.760 13.700 56.400 ;
        RECT 10.900 54.400 11.770 55.760 ;
        RECT 18.850 55.750 19.200 57.400 ;
        RECT 2.800 54.370 3.570 54.400 ;
        RECT 2.800 53.410 3.580 54.370 ;
        RECT 8.900 54.160 11.770 54.400 ;
        RECT 8.900 53.930 16.930 54.160 ;
        RECT 8.900 53.920 16.890 53.930 ;
        RECT 8.900 53.810 16.880 53.920 ;
        RECT 8.900 53.550 16.860 53.810 ;
        RECT 2.800 52.510 3.570 53.410 ;
        RECT 8.900 53.380 16.940 53.550 ;
        RECT 9.600 53.320 16.940 53.380 ;
        RECT 9.600 53.300 13.310 53.320 ;
        RECT 9.600 52.990 12.800 53.300 ;
        RECT 2.800 51.680 3.800 52.510 ;
        RECT 9.600 52.310 11.780 52.990 ;
        RECT 9.600 52.300 11.760 52.310 ;
        RECT 3.170 43.700 3.800 51.680 ;
        RECT 0.790 42.600 4.010 43.700 ;
        RECT 0.800 42.350 1.000 42.600 ;
        RECT 0.790 41.390 1.020 42.350 ;
        RECT 0.800 41.060 1.000 41.390 ;
        RECT 0.790 40.100 1.020 41.060 ;
        RECT 0.800 39.770 1.000 40.100 ;
        RECT 0.790 38.810 1.020 39.770 ;
        RECT 0.800 38.790 1.000 38.810 ;
      LAYER via ;
        RECT 18.300 57.600 18.590 58.200 ;
        RECT 12.800 55.910 13.500 56.200 ;
      LAYER met2 ;
        RECT 18.200 56.300 18.700 58.400 ;
        RECT 12.700 55.800 18.700 56.300 ;
    END
  END Ptatin
  PIN GND
    ANTENNADIFFAREA 7.540000 ;
    PORT
      LAYER li1 ;
        RECT 19.340 61.980 25.380 62.150 ;
        RECT 11.910 55.250 16.950 55.420 ;
        RECT 3.720 53.160 8.760 53.330 ;
        RECT 11.920 52.060 16.960 52.230 ;
        RECT -4.390 38.560 0.650 38.730 ;
      LAYER mcon ;
        RECT 19.420 61.980 25.300 62.150 ;
        RECT 11.990 55.250 16.870 55.420 ;
        RECT 3.800 53.160 8.680 53.330 ;
        RECT 12.000 52.060 16.880 52.230 ;
        RECT -4.310 38.560 0.570 38.730 ;
      LAYER met1 ;
        RECT 14.900 62.330 25.310 62.810 ;
        RECT 14.900 62.300 19.200 62.330 ;
        RECT 19.460 62.320 25.310 62.330 ;
        RECT 14.900 58.500 16.620 62.300 ;
        RECT 19.460 62.180 25.240 62.320 ;
        RECT 19.360 61.950 25.360 62.180 ;
        RECT 14.800 56.400 15.700 57.510 ;
        RECT 14.800 56.100 17.500 56.400 ;
        RECT 17.100 55.510 17.500 56.100 ;
        RECT 11.990 55.450 17.500 55.510 ;
        RECT 11.930 55.240 17.500 55.450 ;
        RECT 11.930 55.220 16.930 55.240 ;
        RECT 3.750 53.360 8.720 53.370 ;
        RECT 3.740 53.130 8.740 53.360 ;
        RECT 3.750 53.010 8.720 53.130 ;
        RECT 7.200 51.500 8.690 53.010 ;
        RECT 17.100 52.270 17.500 55.240 ;
        RECT 12.000 52.260 17.500 52.270 ;
        RECT 11.940 52.030 17.500 52.260 ;
        RECT 12.000 52.000 17.500 52.030 ;
        RECT 17.100 51.510 17.500 52.000 ;
        RECT 16.190 51.500 17.500 51.510 ;
        RECT 7.200 50.800 17.500 51.500 ;
        RECT -4.370 38.700 0.630 38.760 ;
        RECT 16.190 38.700 17.500 50.800 ;
        RECT -4.370 38.650 0.650 38.700 ;
        RECT 1.200 38.650 19.700 38.700 ;
        RECT -4.370 38.530 19.700 38.650 ;
        RECT -4.300 38.100 19.700 38.530 ;
      LAYER via ;
        RECT 15.000 58.600 15.600 58.900 ;
        RECT 15.000 57.000 15.400 57.400 ;
      LAYER met2 ;
        RECT 14.900 56.900 15.700 59.010 ;
    END
  END GND
  PIN Vout
    ANTENNADIFFAREA 3.770000 ;
    PORT
      LAYER li1 ;
        RECT 19.340 55.530 25.380 55.700 ;
        RECT 18.630 52.700 19.670 52.870 ;
        RECT 26.790 26.850 32.830 27.020 ;
      LAYER mcon ;
        RECT 19.420 55.530 25.300 55.700 ;
        RECT 18.710 52.700 19.590 52.870 ;
        RECT 26.870 26.850 32.750 27.020 ;
      LAYER met1 ;
        RECT 19.360 55.500 25.360 55.730 ;
        RECT 20.100 54.800 25.300 55.500 ;
        RECT 18.650 52.900 19.600 52.910 ;
        RECT 18.650 52.750 19.650 52.900 ;
        RECT 18.600 52.670 19.650 52.750 ;
        RECT 18.600 52.160 19.600 52.670 ;
        RECT 22.290 26.860 25.610 28.310 ;
        RECT 26.810 27.020 32.810 27.050 ;
        RECT 26.770 26.860 32.820 27.020 ;
        RECT 22.290 26.500 32.820 26.860 ;
        RECT 22.290 26.490 25.610 26.500 ;
      LAYER via ;
        RECT 22.580 54.900 23.100 55.200 ;
        RECT 18.800 52.200 19.300 52.500 ;
        RECT 23.890 27.310 25.490 28.200 ;
      LAYER met2 ;
        RECT 18.700 52.000 19.360 52.530 ;
        RECT 18.500 51.500 19.510 52.000 ;
        RECT 22.400 30.000 23.300 55.400 ;
        RECT 22.400 27.850 25.910 30.000 ;
        RECT 23.770 27.190 25.910 27.850 ;
      LAYER via2 ;
        RECT 18.800 51.600 19.300 51.900 ;
        RECT 23.800 28.410 25.500 28.700 ;
      LAYER met3 ;
        RECT 7.200 51.510 8.690 53.350 ;
        RECT 18.500 51.510 19.510 52.000 ;
        RECT 2.700 28.310 26.395 51.510 ;
        RECT 23.280 27.850 25.910 28.310 ;
        RECT 23.770 27.190 25.910 27.850 ;
      LAYER via3 ;
        RECT 2.800 28.450 3.120 51.370 ;
      LAYER met4 ;
        RECT 2.720 28.370 3.200 51.450 ;
    END
  END Vout
  PIN VDD
    ANTENNADIFFAREA 7.250000 ;
    PORT
      LAYER li1 ;
        RECT 26.790 62.250 32.830 62.420 ;
        RECT -12.810 61.980 -6.770 62.150 ;
        RECT -4.520 61.980 1.520 62.150 ;
        RECT 3.670 61.930 9.710 62.100 ;
        RECT 11.770 61.890 12.810 62.060 ;
      LAYER mcon ;
        RECT 26.870 62.250 32.750 62.420 ;
        RECT -12.730 61.980 -6.850 62.150 ;
        RECT -4.440 61.980 1.440 62.150 ;
        RECT 3.750 61.930 9.630 62.100 ;
        RECT 11.850 61.890 12.730 62.060 ;
      LAYER met1 ;
        RECT -12.840 63.000 33.000 64.000 ;
        RECT -12.840 61.960 -6.780 63.000 ;
        RECT -4.510 61.970 1.550 63.000 ;
        RECT -12.790 61.950 -6.790 61.960 ;
        RECT -4.500 61.950 1.500 61.970 ;
        RECT 3.690 61.920 9.750 63.000 ;
        RECT 11.840 62.090 12.810 63.000 ;
        RECT 26.830 62.450 33.000 63.000 ;
        RECT 26.810 62.240 33.000 62.450 ;
        RECT 26.810 62.220 32.810 62.240 ;
        RECT 3.690 61.900 9.690 61.920 ;
        RECT 11.790 61.870 12.810 62.090 ;
        RECT 11.790 61.860 12.790 61.870 ;
    END
  END VDD
  OBS
      LAYER nwell ;
        RECT -13.100 48.840 -6.290 62.390 ;
        RECT -5.000 48.840 1.810 62.390 ;
        RECT 3.190 55.240 10.000 62.340 ;
        RECT 11.290 61.210 13.100 62.300 ;
        RECT 11.300 58.800 13.110 59.890 ;
        RECT 11.290 56.390 13.100 57.480 ;
        RECT 26.310 26.610 33.120 62.660 ;
      LAYER li1 ;
        RECT -6.555 60.920 -6.385 61.920 ;
        RECT -4.905 60.920 -4.735 61.920 ;
        RECT 3.285 60.870 3.455 61.870 ;
        RECT 11.385 61.590 11.555 61.920 ;
        RECT 26.405 61.875 26.575 62.205 ;
        RECT 26.790 61.660 32.830 61.830 ;
        RECT 11.770 61.450 12.810 61.620 ;
        RECT 26.405 61.285 26.575 61.615 ;
        RECT 26.790 61.070 32.830 61.240 ;
        RECT -12.810 60.690 -6.770 60.860 ;
        RECT -4.520 60.690 1.520 60.860 ;
        RECT 3.670 60.640 9.710 60.810 ;
        RECT 19.340 60.690 25.380 60.860 ;
        RECT 26.405 60.695 26.575 61.025 ;
        RECT -6.555 59.630 -6.385 60.630 ;
        RECT -4.905 59.630 -4.735 60.630 ;
        RECT 3.285 59.580 3.455 60.580 ;
        RECT 26.790 60.480 32.830 60.650 ;
        RECT 26.405 60.105 26.575 60.435 ;
        RECT 26.790 59.890 32.830 60.060 ;
        RECT -12.810 59.400 -6.770 59.570 ;
        RECT -4.520 59.400 1.520 59.570 ;
        RECT 3.670 59.350 9.710 59.520 ;
        RECT -6.555 58.340 -6.385 59.340 ;
        RECT -4.905 58.340 -4.735 59.340 ;
        RECT 3.285 58.290 3.455 59.290 ;
        RECT 11.395 59.180 11.565 59.510 ;
        RECT 11.780 59.480 12.820 59.650 ;
        RECT 19.340 59.400 25.380 59.570 ;
        RECT 26.405 59.515 26.575 59.845 ;
        RECT 26.790 59.300 32.830 59.470 ;
        RECT 11.780 59.040 12.820 59.210 ;
        RECT 26.405 58.925 26.575 59.255 ;
        RECT 26.790 58.710 32.830 58.880 ;
        RECT 26.405 58.335 26.575 58.665 ;
        RECT -12.810 58.110 -6.770 58.280 ;
        RECT -4.520 58.110 1.520 58.280 ;
        RECT 3.670 58.060 9.710 58.230 ;
        RECT 19.340 58.110 25.380 58.280 ;
        RECT 26.790 58.120 32.830 58.290 ;
        RECT -6.555 57.050 -6.385 58.050 ;
        RECT -4.905 57.050 -4.735 58.050 ;
        RECT 3.285 57.000 3.455 58.000 ;
        RECT 26.405 57.745 26.575 58.075 ;
        RECT 26.790 57.530 32.830 57.700 ;
        RECT 11.770 57.070 12.810 57.240 ;
        RECT 26.405 57.155 26.575 57.485 ;
        RECT -12.810 56.820 -6.770 56.990 ;
        RECT -4.520 56.820 1.520 56.990 ;
        RECT 3.670 56.770 9.710 56.940 ;
        RECT 19.340 56.820 25.380 56.990 ;
        RECT 26.790 56.940 32.830 57.110 ;
        RECT -6.555 55.760 -6.385 56.760 ;
        RECT -4.905 55.760 -4.735 56.760 ;
        RECT 3.285 55.710 3.455 56.710 ;
        RECT 26.405 56.565 26.575 56.895 ;
        RECT 26.790 56.350 32.830 56.520 ;
        RECT 26.405 55.975 26.575 56.305 ;
        RECT 26.790 55.760 32.830 55.930 ;
        RECT -12.810 55.530 -6.770 55.700 ;
        RECT -4.520 55.530 1.520 55.700 ;
        RECT 3.670 55.480 9.710 55.650 ;
        RECT -6.555 54.470 -6.385 55.470 ;
        RECT -4.905 54.470 -4.735 55.470 ;
        RECT 26.405 55.385 26.575 55.715 ;
        RECT 26.790 55.170 32.830 55.340 ;
        RECT 26.405 54.795 26.575 55.125 ;
        RECT 3.720 54.450 8.760 54.620 ;
        RECT 26.790 54.580 32.830 54.750 ;
        RECT -12.810 54.240 -6.770 54.410 ;
        RECT -4.520 54.240 1.520 54.410 ;
        RECT 26.405 54.205 26.575 54.535 ;
        RECT -6.555 53.180 -6.385 54.180 ;
        RECT -4.905 53.180 -4.735 54.180 ;
        RECT 18.630 53.990 19.670 54.160 ;
        RECT 26.790 53.990 32.830 54.160 ;
        RECT -12.810 52.950 -6.770 53.120 ;
        RECT -4.520 52.950 1.520 53.120 ;
        RECT 18.290 52.930 18.460 53.930 ;
        RECT 26.405 53.615 26.575 53.945 ;
        RECT 26.790 53.400 32.830 53.570 ;
        RECT 26.405 53.025 26.575 53.355 ;
        RECT -6.555 51.890 -6.385 52.890 ;
        RECT -4.905 51.890 -4.735 52.890 ;
        RECT 26.790 52.810 32.830 52.980 ;
        RECT 26.405 52.435 26.575 52.765 ;
        RECT 26.790 52.220 32.830 52.390 ;
        RECT 26.405 51.845 26.575 52.175 ;
        RECT -12.810 51.660 -6.770 51.830 ;
        RECT -4.520 51.660 1.520 51.830 ;
        RECT 26.790 51.630 32.830 51.800 ;
        RECT -6.555 50.600 -6.385 51.600 ;
        RECT -4.905 50.600 -4.735 51.600 ;
        RECT 26.405 51.255 26.575 51.585 ;
        RECT 26.790 51.040 32.830 51.210 ;
        RECT 26.405 50.665 26.575 50.995 ;
        RECT -12.810 50.370 -6.770 50.540 ;
        RECT -4.520 50.370 1.520 50.540 ;
        RECT 26.790 50.450 32.830 50.620 ;
        RECT -6.555 49.310 -6.385 50.310 ;
        RECT -4.905 49.310 -4.735 50.310 ;
        RECT 26.405 50.075 26.575 50.405 ;
        RECT 26.790 49.860 32.830 50.030 ;
        RECT 26.405 49.485 26.575 49.815 ;
        RECT 26.790 49.270 32.830 49.440 ;
        RECT -12.810 49.080 -6.770 49.250 ;
        RECT -4.520 49.080 1.520 49.250 ;
        RECT 26.405 48.895 26.575 49.225 ;
        RECT 26.790 48.680 32.830 48.850 ;
        RECT -12.180 48.230 -6.470 48.400 ;
        RECT -4.890 48.230 0.820 48.400 ;
        RECT 26.405 48.305 26.575 48.635 ;
        RECT 26.790 48.090 32.830 48.260 ;
        RECT 26.405 47.715 26.575 48.045 ;
        RECT 26.790 47.500 32.830 47.670 ;
        RECT 26.405 47.125 26.575 47.455 ;
        RECT -12.180 46.940 -6.470 47.110 ;
        RECT -4.890 46.940 0.820 47.110 ;
        RECT 26.790 46.910 32.830 47.080 ;
        RECT 26.405 46.535 26.575 46.865 ;
        RECT 26.790 46.320 32.830 46.490 ;
        RECT 26.405 45.945 26.575 46.275 ;
        RECT -12.180 45.650 -6.470 45.820 ;
        RECT -4.890 45.650 0.820 45.820 ;
        RECT 26.790 45.730 32.830 45.900 ;
        RECT 26.405 45.355 26.575 45.685 ;
        RECT 26.790 45.140 32.830 45.310 ;
        RECT 26.405 44.765 26.575 45.095 ;
        RECT 26.790 44.550 32.830 44.720 ;
        RECT -12.180 44.360 -6.470 44.530 ;
        RECT -4.890 44.360 0.820 44.530 ;
        RECT 26.405 44.175 26.575 44.505 ;
        RECT 26.790 43.960 32.830 44.130 ;
        RECT -4.390 43.720 0.650 43.890 ;
        RECT 26.405 43.585 26.575 43.915 ;
        RECT 26.790 43.370 32.830 43.540 ;
        RECT 26.405 42.995 26.575 43.325 ;
        RECT 26.790 42.780 32.830 42.950 ;
        RECT -4.390 42.430 0.650 42.600 ;
        RECT 26.405 42.405 26.575 42.735 ;
        RECT 26.790 42.190 32.830 42.360 ;
        RECT 26.405 41.815 26.575 42.145 ;
        RECT 26.790 41.600 32.830 41.770 ;
        RECT -4.390 41.140 0.650 41.310 ;
        RECT 26.405 41.225 26.575 41.555 ;
        RECT 26.790 41.010 32.830 41.180 ;
        RECT 26.405 40.635 26.575 40.965 ;
        RECT 26.790 40.420 32.830 40.590 ;
        RECT 26.405 40.045 26.575 40.375 ;
        RECT -4.390 39.850 0.650 40.020 ;
        RECT 26.790 39.830 32.830 40.000 ;
        RECT 26.405 39.455 26.575 39.785 ;
        RECT 26.790 39.240 32.830 39.410 ;
        RECT 26.405 38.865 26.575 39.195 ;
        RECT 26.790 38.650 32.830 38.820 ;
        RECT 26.405 38.275 26.575 38.605 ;
        RECT 26.790 38.060 32.830 38.230 ;
        RECT 26.405 37.685 26.575 38.015 ;
        RECT 26.790 37.470 32.830 37.640 ;
        RECT 26.405 37.095 26.575 37.425 ;
        RECT 26.790 36.880 32.830 37.050 ;
        RECT 26.405 36.505 26.575 36.835 ;
        RECT 26.790 36.290 32.830 36.460 ;
        RECT 26.405 35.915 26.575 36.245 ;
        RECT 26.790 35.700 32.830 35.870 ;
        RECT 26.405 35.325 26.575 35.655 ;
        RECT 26.790 35.110 32.830 35.280 ;
        RECT 26.405 34.735 26.575 35.065 ;
        RECT 26.790 34.520 32.830 34.690 ;
        RECT 26.405 34.145 26.575 34.475 ;
        RECT 26.790 33.930 32.830 34.100 ;
        RECT 26.405 33.555 26.575 33.885 ;
        RECT 26.790 33.340 32.830 33.510 ;
        RECT 26.405 32.965 26.575 33.295 ;
        RECT 26.790 32.750 32.830 32.920 ;
        RECT 26.405 32.375 26.575 32.705 ;
        RECT 26.790 32.160 32.830 32.330 ;
        RECT 26.405 31.785 26.575 32.115 ;
        RECT 26.790 31.570 32.830 31.740 ;
        RECT 26.405 31.195 26.575 31.525 ;
        RECT 26.790 30.980 32.830 31.150 ;
        RECT 26.405 30.605 26.575 30.935 ;
        RECT 26.790 30.390 32.830 30.560 ;
        RECT 26.405 30.015 26.575 30.345 ;
        RECT 26.790 29.800 32.830 29.970 ;
        RECT 26.405 29.425 26.575 29.755 ;
        RECT 26.790 29.210 32.830 29.380 ;
        RECT 26.405 28.835 26.575 29.165 ;
        RECT 26.790 28.620 32.830 28.790 ;
        RECT 26.405 28.245 26.575 28.575 ;
        RECT 26.790 28.030 32.830 28.200 ;
        RECT 26.405 27.655 26.575 27.985 ;
        RECT 26.790 27.440 32.830 27.610 ;
        RECT 26.405 27.065 26.575 27.395 ;
      LAYER mcon ;
        RECT 26.405 61.955 26.575 62.125 ;
        RECT -6.555 61.000 -6.385 61.840 ;
        RECT -4.905 61.000 -4.735 61.840 ;
        RECT 3.285 60.950 3.455 61.790 ;
        RECT 11.385 61.670 11.555 61.840 ;
        RECT 26.870 61.660 32.750 61.830 ;
        RECT 11.850 61.450 12.730 61.620 ;
        RECT 26.405 61.365 26.575 61.535 ;
        RECT 26.870 61.070 32.750 61.240 ;
        RECT -12.730 60.690 -6.850 60.860 ;
        RECT -4.440 60.690 1.440 60.860 ;
        RECT 3.750 60.640 9.630 60.810 ;
        RECT 19.420 60.690 25.300 60.860 ;
        RECT 26.405 60.775 26.575 60.945 ;
        RECT -6.555 59.710 -6.385 60.550 ;
        RECT -4.905 59.710 -4.735 60.550 ;
        RECT 3.285 59.660 3.455 60.500 ;
        RECT 26.870 60.480 32.750 60.650 ;
        RECT 26.405 60.185 26.575 60.355 ;
        RECT 26.870 59.890 32.750 60.060 ;
        RECT -12.730 59.400 -6.850 59.570 ;
        RECT -4.440 59.400 1.440 59.570 ;
        RECT 3.750 59.350 9.630 59.520 ;
        RECT 11.860 59.480 12.740 59.650 ;
        RECT 26.405 59.595 26.575 59.765 ;
        RECT -6.555 58.420 -6.385 59.260 ;
        RECT -4.905 58.420 -4.735 59.260 ;
        RECT 3.285 58.370 3.455 59.210 ;
        RECT 11.395 59.260 11.565 59.430 ;
        RECT 19.420 59.400 25.300 59.570 ;
        RECT 26.870 59.300 32.750 59.470 ;
        RECT 11.860 59.040 12.740 59.210 ;
        RECT 26.405 59.005 26.575 59.175 ;
        RECT 26.870 58.710 32.750 58.880 ;
        RECT 26.405 58.415 26.575 58.585 ;
        RECT -12.730 58.110 -6.850 58.280 ;
        RECT -4.440 58.110 1.440 58.280 ;
        RECT 3.750 58.060 9.630 58.230 ;
        RECT 19.420 58.110 25.300 58.280 ;
        RECT 26.870 58.120 32.750 58.290 ;
        RECT -6.555 57.130 -6.385 57.970 ;
        RECT -4.905 57.130 -4.735 57.970 ;
        RECT 3.285 57.080 3.455 57.920 ;
        RECT 26.405 57.825 26.575 57.995 ;
        RECT 26.870 57.530 32.750 57.700 ;
        RECT 11.850 57.070 12.730 57.240 ;
        RECT 26.405 57.235 26.575 57.405 ;
        RECT -12.730 56.820 -6.850 56.990 ;
        RECT -4.440 56.820 1.440 56.990 ;
        RECT 3.750 56.770 9.630 56.940 ;
        RECT 19.420 56.820 25.300 56.990 ;
        RECT 26.870 56.940 32.750 57.110 ;
        RECT -6.555 55.840 -6.385 56.680 ;
        RECT -4.905 55.840 -4.735 56.680 ;
        RECT 3.285 55.790 3.455 56.630 ;
        RECT 26.405 56.645 26.575 56.815 ;
        RECT 26.870 56.350 32.750 56.520 ;
        RECT 26.405 56.055 26.575 56.225 ;
        RECT 26.870 55.760 32.750 55.930 ;
        RECT -12.730 55.530 -6.850 55.700 ;
        RECT -4.440 55.530 1.440 55.700 ;
        RECT 3.750 55.480 9.630 55.650 ;
        RECT -6.555 54.550 -6.385 55.390 ;
        RECT -4.905 54.550 -4.735 55.390 ;
        RECT 26.405 55.465 26.575 55.635 ;
        RECT 26.870 55.170 32.750 55.340 ;
        RECT 26.405 54.875 26.575 55.045 ;
        RECT 3.800 54.450 8.680 54.620 ;
        RECT 26.870 54.580 32.750 54.750 ;
        RECT -12.730 54.240 -6.850 54.410 ;
        RECT -4.440 54.240 1.440 54.410 ;
        RECT 26.405 54.285 26.575 54.455 ;
        RECT -6.555 53.260 -6.385 54.100 ;
        RECT -4.905 53.260 -4.735 54.100 ;
        RECT 18.710 53.990 19.590 54.160 ;
        RECT 26.870 53.990 32.750 54.160 ;
        RECT -12.730 52.950 -6.850 53.120 ;
        RECT -4.440 52.950 1.440 53.120 ;
        RECT 18.290 53.010 18.460 53.850 ;
        RECT 26.405 53.695 26.575 53.865 ;
        RECT 26.870 53.400 32.750 53.570 ;
        RECT 26.405 53.105 26.575 53.275 ;
        RECT -6.555 51.970 -6.385 52.810 ;
        RECT 26.870 52.810 32.750 52.980 ;
        RECT -4.905 51.970 -4.735 52.810 ;
        RECT 26.405 52.515 26.575 52.685 ;
        RECT 26.870 52.220 32.750 52.390 ;
        RECT 26.405 51.925 26.575 52.095 ;
        RECT -12.730 51.660 -6.850 51.830 ;
        RECT -4.440 51.660 1.440 51.830 ;
        RECT 26.870 51.630 32.750 51.800 ;
        RECT -6.555 50.680 -6.385 51.520 ;
        RECT -4.905 50.680 -4.735 51.520 ;
        RECT 26.405 51.335 26.575 51.505 ;
        RECT 26.870 51.040 32.750 51.210 ;
        RECT 26.405 50.745 26.575 50.915 ;
        RECT -12.730 50.370 -6.850 50.540 ;
        RECT -4.440 50.370 1.440 50.540 ;
        RECT 26.870 50.450 32.750 50.620 ;
        RECT -6.555 49.390 -6.385 50.230 ;
        RECT -4.905 49.390 -4.735 50.230 ;
        RECT 26.405 50.155 26.575 50.325 ;
        RECT 26.870 49.860 32.750 50.030 ;
        RECT 26.405 49.565 26.575 49.735 ;
        RECT 26.870 49.270 32.750 49.440 ;
        RECT -12.730 49.080 -6.850 49.250 ;
        RECT -4.440 49.080 1.440 49.250 ;
        RECT 26.405 48.975 26.575 49.145 ;
        RECT 26.870 48.680 32.750 48.850 ;
        RECT -12.100 48.230 -6.550 48.400 ;
        RECT -4.810 48.230 0.740 48.400 ;
        RECT 26.405 48.385 26.575 48.555 ;
        RECT 26.870 48.090 32.750 48.260 ;
        RECT 26.405 47.795 26.575 47.965 ;
        RECT 26.870 47.500 32.750 47.670 ;
        RECT 26.405 47.205 26.575 47.375 ;
        RECT -12.100 46.940 -6.550 47.110 ;
        RECT -4.810 46.940 0.740 47.110 ;
        RECT 26.870 46.910 32.750 47.080 ;
        RECT 26.405 46.615 26.575 46.785 ;
        RECT 26.870 46.320 32.750 46.490 ;
        RECT 26.405 46.025 26.575 46.195 ;
        RECT -12.100 45.650 -6.550 45.820 ;
        RECT -4.810 45.650 0.740 45.820 ;
        RECT 26.870 45.730 32.750 45.900 ;
        RECT 26.405 45.435 26.575 45.605 ;
        RECT 26.870 45.140 32.750 45.310 ;
        RECT 26.405 44.845 26.575 45.015 ;
        RECT 26.870 44.550 32.750 44.720 ;
        RECT -12.100 44.360 -6.550 44.530 ;
        RECT -4.810 44.360 0.740 44.530 ;
        RECT 26.405 44.255 26.575 44.425 ;
        RECT 26.870 43.960 32.750 44.130 ;
        RECT -4.310 43.720 0.570 43.890 ;
        RECT 26.405 43.665 26.575 43.835 ;
        RECT 26.870 43.370 32.750 43.540 ;
        RECT 26.405 43.075 26.575 43.245 ;
        RECT 26.870 42.780 32.750 42.950 ;
        RECT -4.310 42.430 0.570 42.600 ;
        RECT 26.405 42.485 26.575 42.655 ;
        RECT 26.870 42.190 32.750 42.360 ;
        RECT 26.405 41.895 26.575 42.065 ;
        RECT 26.870 41.600 32.750 41.770 ;
        RECT -4.310 41.140 0.570 41.310 ;
        RECT 26.405 41.305 26.575 41.475 ;
        RECT 26.870 41.010 32.750 41.180 ;
        RECT 26.405 40.715 26.575 40.885 ;
        RECT 26.870 40.420 32.750 40.590 ;
        RECT 26.405 40.125 26.575 40.295 ;
        RECT -4.310 39.850 0.570 40.020 ;
        RECT 26.870 39.830 32.750 40.000 ;
        RECT 26.405 39.535 26.575 39.705 ;
        RECT 26.870 39.240 32.750 39.410 ;
        RECT 26.405 38.945 26.575 39.115 ;
        RECT 26.870 38.650 32.750 38.820 ;
        RECT 26.405 38.355 26.575 38.525 ;
        RECT 26.870 38.060 32.750 38.230 ;
        RECT 26.405 37.765 26.575 37.935 ;
        RECT 26.870 37.470 32.750 37.640 ;
        RECT 26.405 37.175 26.575 37.345 ;
        RECT 26.870 36.880 32.750 37.050 ;
        RECT 26.405 36.585 26.575 36.755 ;
        RECT 26.870 36.290 32.750 36.460 ;
        RECT 26.405 35.995 26.575 36.165 ;
        RECT 26.870 35.700 32.750 35.870 ;
        RECT 26.405 35.405 26.575 35.575 ;
        RECT 26.870 35.110 32.750 35.280 ;
        RECT 26.405 34.815 26.575 34.985 ;
        RECT 26.870 34.520 32.750 34.690 ;
        RECT 26.405 34.225 26.575 34.395 ;
        RECT 26.870 33.930 32.750 34.100 ;
        RECT 26.405 33.635 26.575 33.805 ;
        RECT 26.870 33.340 32.750 33.510 ;
        RECT 26.405 33.045 26.575 33.215 ;
        RECT 26.870 32.750 32.750 32.920 ;
        RECT 26.405 32.455 26.575 32.625 ;
        RECT 26.870 32.160 32.750 32.330 ;
        RECT 26.405 31.865 26.575 32.035 ;
        RECT 26.870 31.570 32.750 31.740 ;
        RECT 26.405 31.275 26.575 31.445 ;
        RECT 26.870 30.980 32.750 31.150 ;
        RECT 26.405 30.685 26.575 30.855 ;
        RECT 26.870 30.390 32.750 30.560 ;
        RECT 26.405 30.095 26.575 30.265 ;
        RECT 26.870 29.800 32.750 29.970 ;
        RECT 26.405 29.505 26.575 29.675 ;
        RECT 26.870 29.210 32.750 29.380 ;
        RECT 26.405 28.915 26.575 29.085 ;
        RECT 26.870 28.620 32.750 28.790 ;
        RECT 26.405 28.325 26.575 28.495 ;
        RECT 26.870 28.030 32.750 28.200 ;
        RECT 26.405 27.735 26.575 27.905 ;
        RECT 26.870 27.440 32.750 27.610 ;
        RECT 26.405 27.145 26.575 27.315 ;
      LAYER met1 ;
        RECT 26.300 62.185 26.600 62.200 ;
        RECT -12.790 60.660 -6.790 60.890 ;
        RECT -12.790 59.370 -6.790 59.600 ;
        RECT -12.790 58.080 -6.790 58.310 ;
        RECT -12.790 56.790 -6.790 57.020 ;
        RECT -12.790 55.500 -6.790 55.730 ;
        RECT -12.790 54.210 -6.790 54.440 ;
        RECT -12.790 52.920 -6.790 53.150 ;
        RECT -12.790 51.630 -6.790 51.860 ;
        RECT -12.790 50.340 -6.790 50.570 ;
        RECT -6.600 49.300 -4.700 61.900 ;
        RECT -4.500 60.660 1.500 60.890 ;
        RECT 3.200 60.600 3.500 61.900 ;
        RECT 11.300 61.200 11.630 61.910 ;
        RECT 26.300 61.895 26.605 62.185 ;
        RECT 11.790 61.620 12.790 61.650 ;
        RECT 11.790 61.420 12.800 61.620 ;
        RECT 11.800 61.200 12.800 61.420 ;
        RECT 11.300 61.000 12.800 61.200 ;
        RECT 3.690 60.610 9.690 60.840 ;
        RECT -4.500 59.370 1.500 59.600 ;
        RECT 2.200 59.300 3.500 60.600 ;
        RECT 3.690 59.320 9.690 59.550 ;
        RECT -4.500 58.080 1.500 58.310 ;
        RECT -4.500 56.790 1.500 57.020 ;
        RECT -4.500 55.500 1.500 55.730 ;
        RECT 3.200 55.700 3.500 59.300 ;
        RECT 11.290 58.800 11.620 59.510 ;
        RECT 11.800 59.450 12.800 61.000 ;
        RECT 26.300 61.595 26.600 61.895 ;
        RECT 26.810 61.630 32.810 61.860 ;
        RECT 26.300 61.305 26.605 61.595 ;
        RECT 26.300 61.005 26.600 61.305 ;
        RECT 26.810 61.040 32.810 61.270 ;
        RECT 19.360 60.660 25.360 60.890 ;
        RECT 26.300 60.715 26.605 61.005 ;
        RECT 26.300 60.415 26.600 60.715 ;
        RECT 26.810 60.450 32.810 60.680 ;
        RECT 26.300 60.125 26.605 60.415 ;
        RECT 26.300 59.825 26.600 60.125 ;
        RECT 26.810 59.860 32.810 60.090 ;
        RECT 19.360 59.370 25.360 59.600 ;
        RECT 26.300 59.535 26.605 59.825 ;
        RECT 11.800 58.800 12.800 59.240 ;
        RECT 11.290 58.600 12.800 58.800 ;
        RECT 3.690 58.030 9.690 58.260 ;
        RECT 11.800 58.110 12.800 58.600 ;
        RECT 26.300 59.235 26.600 59.535 ;
        RECT 26.810 59.270 32.810 59.500 ;
        RECT 26.300 58.945 26.605 59.235 ;
        RECT 26.300 58.645 26.600 58.945 ;
        RECT 26.810 58.680 32.810 58.910 ;
        RECT 26.300 58.355 26.605 58.645 ;
        RECT 11.800 57.700 17.700 58.110 ;
        RECT 19.360 58.080 25.360 58.310 ;
        RECT 11.800 57.270 12.800 57.700 ;
        RECT 11.790 57.070 12.800 57.270 ;
        RECT 17.200 57.100 17.700 57.700 ;
        RECT 26.300 58.055 26.600 58.355 ;
        RECT 26.810 58.090 32.810 58.320 ;
        RECT 26.300 57.765 26.605 58.055 ;
        RECT 26.300 57.465 26.600 57.765 ;
        RECT 26.810 57.500 32.810 57.730 ;
        RECT 26.300 57.175 26.605 57.465 ;
        RECT 11.790 57.040 12.790 57.070 ;
        RECT 3.690 56.740 9.690 56.970 ;
        RECT 17.200 56.700 18.080 57.100 ;
        RECT 19.360 56.790 25.360 57.020 ;
        RECT 26.300 56.875 26.600 57.175 ;
        RECT 26.810 56.910 32.810 57.140 ;
        RECT 3.690 55.450 9.690 55.680 ;
        RECT 3.800 54.650 8.700 55.450 ;
        RECT -4.500 54.210 1.500 54.440 ;
        RECT 3.740 54.420 8.740 54.650 ;
        RECT 3.800 54.400 8.700 54.420 ;
        RECT 17.720 53.900 18.080 56.700 ;
        RECT 26.300 56.585 26.605 56.875 ;
        RECT 26.300 56.285 26.600 56.585 ;
        RECT 26.810 56.320 32.810 56.550 ;
        RECT 26.300 55.995 26.605 56.285 ;
        RECT 26.300 55.695 26.600 55.995 ;
        RECT 26.810 55.730 32.810 55.960 ;
        RECT 26.300 55.405 26.605 55.695 ;
        RECT 18.600 54.190 19.620 55.210 ;
        RECT 26.300 55.105 26.600 55.405 ;
        RECT 26.810 55.140 32.810 55.370 ;
        RECT 26.300 54.815 26.605 55.105 ;
        RECT 26.300 54.515 26.600 54.815 ;
        RECT 26.810 54.550 32.810 54.780 ;
        RECT 26.300 54.225 26.605 54.515 ;
        RECT 18.600 54.100 19.650 54.190 ;
        RECT 18.650 53.960 19.650 54.100 ;
        RECT 18.700 53.940 19.620 53.960 ;
        RECT 26.300 53.925 26.600 54.225 ;
        RECT 26.810 53.960 32.810 54.190 ;
        RECT 18.260 53.900 18.490 53.910 ;
        RECT -4.500 52.920 1.500 53.150 ;
        RECT 17.720 52.900 18.500 53.900 ;
        RECT 26.300 53.635 26.605 53.925 ;
        RECT 26.300 53.335 26.600 53.635 ;
        RECT 26.810 53.370 32.810 53.600 ;
        RECT 26.300 53.045 26.605 53.335 ;
        RECT 26.300 52.745 26.600 53.045 ;
        RECT 26.810 52.780 32.810 53.010 ;
        RECT 26.300 52.455 26.605 52.745 ;
        RECT 26.300 52.155 26.600 52.455 ;
        RECT 26.810 52.190 32.810 52.420 ;
        RECT -4.500 51.630 1.500 51.860 ;
        RECT 18.500 51.500 19.510 52.000 ;
        RECT 26.300 51.865 26.605 52.155 ;
        RECT 26.300 51.565 26.600 51.865 ;
        RECT 26.810 51.600 32.810 51.830 ;
        RECT 26.300 51.275 26.605 51.565 ;
        RECT 26.300 50.975 26.600 51.275 ;
        RECT 26.810 51.010 32.810 51.240 ;
        RECT 26.300 50.685 26.605 50.975 ;
        RECT -4.500 50.340 1.500 50.570 ;
        RECT 26.300 50.385 26.600 50.685 ;
        RECT 26.810 50.420 32.810 50.650 ;
        RECT 26.300 50.095 26.605 50.385 ;
        RECT 26.300 49.795 26.600 50.095 ;
        RECT 26.810 49.830 32.810 50.060 ;
        RECT 26.300 49.505 26.605 49.795 ;
        RECT -12.800 49.280 -6.800 49.300 ;
        RECT -12.800 49.050 -6.790 49.280 ;
        RECT -12.800 48.900 -6.800 49.050 ;
        RECT -6.510 48.900 -5.600 49.300 ;
        RECT -12.800 48.400 -5.600 48.900 ;
        RECT -4.510 48.800 1.500 49.300 ;
        RECT 26.300 49.290 26.600 49.505 ;
        RECT -12.160 48.200 -5.600 48.400 ;
        RECT -4.900 48.430 0.300 48.800 ;
        RECT -4.900 48.200 0.800 48.430 ;
        RECT 20.100 48.410 26.610 49.290 ;
        RECT 26.810 49.240 32.810 49.470 ;
        RECT 26.810 48.650 32.810 48.880 ;
        RECT 26.300 48.325 26.605 48.410 ;
        RECT 26.300 48.025 26.600 48.325 ;
        RECT 26.810 48.060 32.810 48.290 ;
        RECT 26.300 47.735 26.605 48.025 ;
        RECT 26.300 47.435 26.600 47.735 ;
        RECT 26.810 47.470 32.810 47.700 ;
        RECT 26.300 47.145 26.605 47.435 ;
        RECT -12.160 46.910 -6.490 47.140 ;
        RECT -4.870 46.910 0.800 47.140 ;
        RECT 26.300 46.845 26.600 47.145 ;
        RECT 26.810 46.880 32.810 47.110 ;
        RECT 26.300 46.555 26.605 46.845 ;
        RECT 26.300 46.255 26.600 46.555 ;
        RECT 26.810 46.290 32.810 46.520 ;
        RECT 26.300 45.965 26.605 46.255 ;
        RECT -12.160 45.620 -6.490 45.850 ;
        RECT -4.870 45.620 0.800 45.850 ;
        RECT 26.300 45.665 26.600 45.965 ;
        RECT 26.810 45.700 32.810 45.930 ;
        RECT 26.300 45.375 26.605 45.665 ;
        RECT 26.300 45.075 26.600 45.375 ;
        RECT 26.810 45.110 32.810 45.340 ;
        RECT 26.300 44.785 26.605 45.075 ;
        RECT -12.160 44.330 0.800 44.560 ;
        RECT 26.300 44.485 26.600 44.785 ;
        RECT 26.810 44.520 32.810 44.750 ;
        RECT -12.120 43.960 0.600 44.330 ;
        RECT -10.760 43.920 0.600 43.960 ;
        RECT 26.300 44.195 26.605 44.485 ;
        RECT -10.760 43.900 0.630 43.920 ;
        RECT -4.690 43.890 0.630 43.900 ;
        RECT -4.370 43.690 0.630 43.890 ;
        RECT 26.300 43.895 26.600 44.195 ;
        RECT 26.810 43.930 32.810 44.160 ;
        RECT 26.300 43.605 26.605 43.895 ;
        RECT 26.300 43.305 26.600 43.605 ;
        RECT 26.810 43.340 32.810 43.570 ;
        RECT 26.300 43.015 26.605 43.305 ;
        RECT 26.300 42.715 26.600 43.015 ;
        RECT 26.810 42.750 32.810 42.980 ;
        RECT -4.370 42.400 0.630 42.630 ;
        RECT 26.300 42.425 26.605 42.715 ;
        RECT 26.300 42.125 26.600 42.425 ;
        RECT 26.810 42.160 32.810 42.390 ;
        RECT 26.300 41.835 26.605 42.125 ;
        RECT 26.300 41.535 26.600 41.835 ;
        RECT 26.810 41.570 32.810 41.800 ;
        RECT -4.370 41.110 0.630 41.340 ;
        RECT 26.300 41.245 26.605 41.535 ;
        RECT 26.300 40.945 26.600 41.245 ;
        RECT 26.810 40.980 32.810 41.210 ;
        RECT 26.300 40.655 26.605 40.945 ;
        RECT 26.300 40.355 26.600 40.655 ;
        RECT 26.810 40.390 32.810 40.620 ;
        RECT 26.300 40.065 26.605 40.355 ;
        RECT -4.370 39.820 0.630 40.050 ;
        RECT 26.300 39.765 26.600 40.065 ;
        RECT 26.810 39.800 32.810 40.030 ;
        RECT 26.300 39.475 26.605 39.765 ;
        RECT 26.300 39.175 26.600 39.475 ;
        RECT 26.810 39.210 32.810 39.440 ;
        RECT 26.300 38.885 26.605 39.175 ;
        RECT 26.300 38.585 26.600 38.885 ;
        RECT 26.810 38.620 32.810 38.850 ;
        RECT 26.300 38.295 26.605 38.585 ;
        RECT 26.300 37.995 26.600 38.295 ;
        RECT 26.810 38.030 32.810 38.260 ;
        RECT 26.300 37.705 26.605 37.995 ;
        RECT 26.300 37.405 26.600 37.705 ;
        RECT 26.810 37.440 32.810 37.670 ;
        RECT 26.300 37.115 26.605 37.405 ;
        RECT 26.300 36.815 26.600 37.115 ;
        RECT 26.810 36.850 32.810 37.080 ;
        RECT 26.300 36.525 26.605 36.815 ;
        RECT 26.300 36.225 26.600 36.525 ;
        RECT 26.810 36.260 32.810 36.490 ;
        RECT 26.300 35.935 26.605 36.225 ;
        RECT 26.300 35.635 26.600 35.935 ;
        RECT 26.810 35.670 32.810 35.900 ;
        RECT 26.300 35.345 26.605 35.635 ;
        RECT 26.300 35.045 26.600 35.345 ;
        RECT 26.810 35.080 32.810 35.310 ;
        RECT 26.300 34.755 26.605 35.045 ;
        RECT 26.300 34.455 26.600 34.755 ;
        RECT 26.810 34.490 32.810 34.720 ;
        RECT 26.300 34.165 26.605 34.455 ;
        RECT 26.300 33.865 26.600 34.165 ;
        RECT 26.810 33.900 32.810 34.130 ;
        RECT 26.300 33.575 26.605 33.865 ;
        RECT 26.300 33.275 26.600 33.575 ;
        RECT 26.810 33.310 32.810 33.540 ;
        RECT 26.300 32.985 26.605 33.275 ;
        RECT 26.300 32.685 26.600 32.985 ;
        RECT 26.810 32.720 32.810 32.950 ;
        RECT 26.300 32.395 26.605 32.685 ;
        RECT 26.300 32.095 26.600 32.395 ;
        RECT 26.810 32.130 32.810 32.360 ;
        RECT 26.300 31.805 26.605 32.095 ;
        RECT 26.300 31.505 26.600 31.805 ;
        RECT 26.810 31.540 32.810 31.770 ;
        RECT 26.300 31.215 26.605 31.505 ;
        RECT 26.300 30.915 26.600 31.215 ;
        RECT 26.810 30.950 32.810 31.180 ;
        RECT 26.300 30.625 26.605 30.915 ;
        RECT 26.300 30.325 26.600 30.625 ;
        RECT 26.810 30.360 32.810 30.590 ;
        RECT 26.300 30.035 26.605 30.325 ;
        RECT 26.300 29.735 26.600 30.035 ;
        RECT 26.810 29.770 32.810 30.000 ;
        RECT 26.300 29.445 26.605 29.735 ;
        RECT 26.300 29.145 26.600 29.445 ;
        RECT 26.810 29.180 32.810 29.410 ;
        RECT 26.300 28.855 26.605 29.145 ;
        RECT 26.300 28.555 26.600 28.855 ;
        RECT 26.810 28.590 32.810 28.820 ;
        RECT 26.300 28.265 26.605 28.555 ;
        RECT 26.300 27.965 26.600 28.265 ;
        RECT 26.810 28.000 32.810 28.230 ;
        RECT 26.300 27.675 26.605 27.965 ;
        RECT 26.300 27.375 26.600 27.675 ;
        RECT 26.810 27.410 32.810 27.640 ;
        RECT 26.300 27.085 26.605 27.375 ;
        RECT 26.300 27.000 26.600 27.085 ;
      LAYER via ;
        RECT -6.000 59.700 -5.400 60.200 ;
        RECT 2.300 59.700 2.900 60.200 ;
        RECT 5.900 54.800 6.600 55.200 ;
        RECT 18.700 54.800 19.500 55.100 ;
        RECT -1.500 48.500 -0.800 48.800 ;
        RECT 20.200 48.600 20.900 49.100 ;
      LAYER met2 ;
        RECT -6.200 59.500 3.000 60.400 ;
        RECT 5.800 55.200 6.700 55.300 ;
        RECT 5.800 54.700 19.610 55.200 ;
        RECT -1.610 48.410 21.100 49.300 ;
      LAYER met4 ;
        RECT 18.400 50.815 19.600 52.000 ;
        RECT 3.890 29.005 25.700 50.815 ;
  END
END tt_um_mete_opamp
END LIBRARY

