magic
tech sky130B
magscale 1 2
timestamp 1768734963
<< metal3 >>
rect -2370 2292 2369 2320
rect -2370 -2292 2285 2292
rect 2349 -2292 2369 2292
rect -2370 -2320 2369 -2292
<< via3 >>
rect 2285 -2292 2349 2292
<< mimcap >>
rect -2270 2180 2170 2220
rect -2270 -2180 -2230 2180
rect 2130 -2180 2170 2180
rect -2270 -2220 2170 -2180
<< mimcapcontact >>
rect -2230 -2180 2130 2180
<< metal4 >>
rect 2269 2292 2365 2308
rect -2231 2180 2131 2181
rect -2231 -2180 -2230 2180
rect 2130 -2180 2131 2180
rect -2231 -2181 2131 -2180
rect 2269 -2292 2285 2292
rect 2349 -2292 2365 2292
rect 2269 -2308 2365 -2292
<< properties >>
string FIXED_BBOX -2370 -2320 2270 2320
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 22.2 l 22.2 val 1.002k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
