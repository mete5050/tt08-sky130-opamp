magic
tech sky130B
magscale 1 2
timestamp 1768756364
<< nmos >>
rect -487 -531 -287 469
rect -229 -531 -29 469
rect 29 -531 229 469
rect 287 -531 487 469
<< ndiff >>
rect -545 457 -487 469
rect -545 -519 -533 457
rect -499 -519 -487 457
rect -545 -531 -487 -519
rect -287 457 -229 469
rect -287 -519 -275 457
rect -241 -519 -229 457
rect -287 -531 -229 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 229 457 287 469
rect 229 -519 241 457
rect 275 -519 287 457
rect 229 -531 287 -519
rect 487 457 545 469
rect 487 -519 499 457
rect 533 -519 545 457
rect 487 -531 545 -519
<< ndiffc >>
rect -533 -519 -499 457
rect -275 -519 -241 457
rect -17 -519 17 457
rect 241 -519 275 457
rect 499 -519 533 457
<< poly >>
rect -487 541 -287 557
rect -487 507 -471 541
rect -303 507 -287 541
rect -487 469 -287 507
rect -229 541 -29 557
rect -229 507 -213 541
rect -45 507 -29 541
rect -229 469 -29 507
rect 29 541 229 557
rect 29 507 45 541
rect 213 507 229 541
rect 29 469 229 507
rect 287 541 487 557
rect 287 507 303 541
rect 471 507 487 541
rect 287 469 487 507
rect -487 -557 -287 -531
rect -229 -557 -29 -531
rect 29 -557 229 -531
rect 287 -557 487 -531
<< polycont >>
rect -471 507 -303 541
rect -213 507 -45 541
rect 45 507 213 541
rect 303 507 471 541
<< locali >>
rect -487 507 -471 541
rect -303 507 -287 541
rect -229 507 -213 541
rect -45 507 -29 541
rect 29 507 45 541
rect 213 507 229 541
rect 287 507 303 541
rect 471 507 487 541
rect -533 457 -499 473
rect -533 -535 -499 -519
rect -275 457 -241 473
rect -275 -535 -241 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 241 457 275 473
rect 241 -535 275 -519
rect 499 457 533 473
rect 499 -535 533 -519
<< viali >>
rect -471 507 -303 541
rect -213 507 -45 541
rect 45 507 213 541
rect 303 507 471 541
rect -533 -519 -499 457
rect -275 -519 -241 457
rect -17 -519 17 457
rect 241 -519 275 457
rect 499 -519 533 457
<< metal1 >>
rect -483 541 -291 547
rect -483 507 -471 541
rect -303 507 -291 541
rect -483 501 -291 507
rect -225 541 -33 547
rect -225 507 -213 541
rect -45 507 -33 541
rect -225 501 -33 507
rect 33 541 225 547
rect 33 507 45 541
rect 213 507 225 541
rect 33 501 225 507
rect 291 541 483 547
rect 291 507 303 541
rect 471 507 483 541
rect 291 501 483 507
rect -539 457 -493 469
rect -539 -519 -533 457
rect -499 -519 -493 457
rect -539 -531 -493 -519
rect -281 457 -235 469
rect -281 -519 -275 457
rect -241 -519 -235 457
rect -281 -531 -235 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 235 457 281 469
rect 235 -519 241 457
rect 275 -519 281 457
rect 235 -531 281 -519
rect 493 457 539 469
rect 493 -519 499 457
rect 533 -519 539 457
rect 493 -531 539 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
