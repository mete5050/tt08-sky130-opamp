magic
tech sky130B
magscale 1 2
timestamp 1768735447
<< nwell >>
rect -1355 -698 1355 664
<< pmos >>
rect -1261 -636 -1061 564
rect -1003 -636 -803 564
rect -745 -636 -545 564
rect -487 -636 -287 564
rect -229 -636 -29 564
rect 29 -636 229 564
rect 287 -636 487 564
rect 545 -636 745 564
rect 803 -636 1003 564
rect 1061 -636 1261 564
<< pdiff >>
rect -1319 552 -1261 564
rect -1319 -624 -1307 552
rect -1273 -624 -1261 552
rect -1319 -636 -1261 -624
rect -1061 552 -1003 564
rect -1061 -624 -1049 552
rect -1015 -624 -1003 552
rect -1061 -636 -1003 -624
rect -803 552 -745 564
rect -803 -624 -791 552
rect -757 -624 -745 552
rect -803 -636 -745 -624
rect -545 552 -487 564
rect -545 -624 -533 552
rect -499 -624 -487 552
rect -545 -636 -487 -624
rect -287 552 -229 564
rect -287 -624 -275 552
rect -241 -624 -229 552
rect -287 -636 -229 -624
rect -29 552 29 564
rect -29 -624 -17 552
rect 17 -624 29 552
rect -29 -636 29 -624
rect 229 552 287 564
rect 229 -624 241 552
rect 275 -624 287 552
rect 229 -636 287 -624
rect 487 552 545 564
rect 487 -624 499 552
rect 533 -624 545 552
rect 487 -636 545 -624
rect 745 552 803 564
rect 745 -624 757 552
rect 791 -624 803 552
rect 745 -636 803 -624
rect 1003 552 1061 564
rect 1003 -624 1015 552
rect 1049 -624 1061 552
rect 1003 -636 1061 -624
rect 1261 552 1319 564
rect 1261 -624 1273 552
rect 1307 -624 1319 552
rect 1261 -636 1319 -624
<< pdiffc >>
rect -1307 -624 -1273 552
rect -1049 -624 -1015 552
rect -791 -624 -757 552
rect -533 -624 -499 552
rect -275 -624 -241 552
rect -17 -624 17 552
rect 241 -624 275 552
rect 499 -624 533 552
rect 757 -624 791 552
rect 1015 -624 1049 552
rect 1273 -624 1307 552
<< poly >>
rect -1261 645 -1061 661
rect -1261 611 -1245 645
rect -1077 611 -1061 645
rect -1261 564 -1061 611
rect -1003 645 -803 661
rect -1003 611 -987 645
rect -819 611 -803 645
rect -1003 564 -803 611
rect -745 645 -545 661
rect -745 611 -729 645
rect -561 611 -545 645
rect -745 564 -545 611
rect -487 645 -287 661
rect -487 611 -471 645
rect -303 611 -287 645
rect -487 564 -287 611
rect -229 645 -29 661
rect -229 611 -213 645
rect -45 611 -29 645
rect -229 564 -29 611
rect 29 645 229 661
rect 29 611 45 645
rect 213 611 229 645
rect 29 564 229 611
rect 287 645 487 661
rect 287 611 303 645
rect 471 611 487 645
rect 287 564 487 611
rect 545 645 745 661
rect 545 611 561 645
rect 729 611 745 645
rect 545 564 745 611
rect 803 645 1003 661
rect 803 611 819 645
rect 987 611 1003 645
rect 803 564 1003 611
rect 1061 645 1261 661
rect 1061 611 1077 645
rect 1245 611 1261 645
rect 1061 564 1261 611
rect -1261 -662 -1061 -636
rect -1003 -662 -803 -636
rect -745 -662 -545 -636
rect -487 -662 -287 -636
rect -229 -662 -29 -636
rect 29 -662 229 -636
rect 287 -662 487 -636
rect 545 -662 745 -636
rect 803 -662 1003 -636
rect 1061 -662 1261 -636
<< polycont >>
rect -1245 611 -1077 645
rect -987 611 -819 645
rect -729 611 -561 645
rect -471 611 -303 645
rect -213 611 -45 645
rect 45 611 213 645
rect 303 611 471 645
rect 561 611 729 645
rect 819 611 987 645
rect 1077 611 1245 645
<< locali >>
rect -1261 611 -1245 645
rect -1077 611 -1061 645
rect -1003 611 -987 645
rect -819 611 -803 645
rect -745 611 -729 645
rect -561 611 -545 645
rect -487 611 -471 645
rect -303 611 -287 645
rect -229 611 -213 645
rect -45 611 -29 645
rect 29 611 45 645
rect 213 611 229 645
rect 287 611 303 645
rect 471 611 487 645
rect 545 611 561 645
rect 729 611 745 645
rect 803 611 819 645
rect 987 611 1003 645
rect 1061 611 1077 645
rect 1245 611 1261 645
rect -1307 552 -1273 568
rect -1307 -640 -1273 -624
rect -1049 552 -1015 568
rect -1049 -640 -1015 -624
rect -791 552 -757 568
rect -791 -640 -757 -624
rect -533 552 -499 568
rect -533 -640 -499 -624
rect -275 552 -241 568
rect -275 -640 -241 -624
rect -17 552 17 568
rect -17 -640 17 -624
rect 241 552 275 568
rect 241 -640 275 -624
rect 499 552 533 568
rect 499 -640 533 -624
rect 757 552 791 568
rect 757 -640 791 -624
rect 1015 552 1049 568
rect 1015 -640 1049 -624
rect 1273 552 1307 568
rect 1273 -640 1307 -624
<< viali >>
rect -1245 611 -1077 645
rect -987 611 -819 645
rect -729 611 -561 645
rect -471 611 -303 645
rect -213 611 -45 645
rect 45 611 213 645
rect 303 611 471 645
rect 561 611 729 645
rect 819 611 987 645
rect 1077 611 1245 645
rect -1307 -624 -1273 552
rect -1049 -624 -1015 552
rect -791 -624 -757 552
rect -533 -624 -499 552
rect -275 -624 -241 552
rect -17 -624 17 552
rect 241 -624 275 552
rect 499 -624 533 552
rect 757 -624 791 552
rect 1015 -624 1049 552
rect 1273 -624 1307 552
<< metal1 >>
rect -1257 645 -1065 651
rect -1257 611 -1245 645
rect -1077 611 -1065 645
rect -1257 605 -1065 611
rect -999 645 -807 651
rect -999 611 -987 645
rect -819 611 -807 645
rect -999 605 -807 611
rect -741 645 -549 651
rect -741 611 -729 645
rect -561 611 -549 645
rect -741 605 -549 611
rect -483 645 -291 651
rect -483 611 -471 645
rect -303 611 -291 645
rect -483 605 -291 611
rect -225 645 -33 651
rect -225 611 -213 645
rect -45 611 -33 645
rect -225 605 -33 611
rect 33 645 225 651
rect 33 611 45 645
rect 213 611 225 645
rect 33 605 225 611
rect 291 645 483 651
rect 291 611 303 645
rect 471 611 483 645
rect 291 605 483 611
rect 549 645 741 651
rect 549 611 561 645
rect 729 611 741 645
rect 549 605 741 611
rect 807 645 999 651
rect 807 611 819 645
rect 987 611 999 645
rect 807 605 999 611
rect 1065 645 1257 651
rect 1065 611 1077 645
rect 1245 611 1257 645
rect 1065 605 1257 611
rect -1313 552 -1267 564
rect -1313 -624 -1307 552
rect -1273 -624 -1267 552
rect -1313 -636 -1267 -624
rect -1055 552 -1009 564
rect -1055 -624 -1049 552
rect -1015 -624 -1009 552
rect -1055 -636 -1009 -624
rect -797 552 -751 564
rect -797 -624 -791 552
rect -757 -624 -751 552
rect -797 -636 -751 -624
rect -539 552 -493 564
rect -539 -624 -533 552
rect -499 -624 -493 552
rect -539 -636 -493 -624
rect -281 552 -235 564
rect -281 -624 -275 552
rect -241 -624 -235 552
rect -281 -636 -235 -624
rect -23 552 23 564
rect -23 -624 -17 552
rect 17 -624 23 552
rect -23 -636 23 -624
rect 235 552 281 564
rect 235 -624 241 552
rect 275 -624 281 552
rect 235 -636 281 -624
rect 493 552 539 564
rect 493 -624 499 552
rect 533 -624 539 552
rect 493 -636 539 -624
rect 751 552 797 564
rect 751 -624 757 552
rect 791 -624 797 552
rect 751 -636 797 -624
rect 1009 552 1055 564
rect 1009 -624 1015 552
rect 1049 -624 1055 552
rect 1009 -636 1055 -624
rect 1267 552 1313 564
rect 1267 -624 1273 552
rect 1307 -624 1313 552
rect 1267 -636 1313 -624
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
