magic
tech sky130B
magscale 1 2
timestamp 1768765927
<< metal1 >>
rect -2568 12600 6600 12800
rect -2568 12392 -1356 12600
rect -902 12394 310 12600
rect 738 12384 1950 12600
rect -1320 12040 -940 12380
rect 640 12120 700 12380
rect 2260 12240 2326 12382
rect 2368 12374 2562 12600
rect 2980 12466 5062 12562
rect 2980 12460 3840 12466
rect 3892 12464 5062 12466
rect 2360 12240 2560 12324
rect 2260 12200 2560 12240
rect -1320 11940 -1200 12040
rect -1080 11940 -940 12040
rect -1320 9860 -940 11940
rect 440 12040 700 12120
rect 440 11940 460 12040
rect 580 11940 700 12040
rect 440 11860 700 11940
rect 640 11140 700 11860
rect 2258 11760 2324 11902
rect 2360 11896 2560 12200
rect 2360 11760 2560 11842
rect 2258 11720 2560 11760
rect 2360 11622 2560 11720
rect 2980 11780 3324 12460
rect 3892 12430 5048 12464
rect 5366 12448 6600 12600
rect 3892 12420 5060 12430
rect 3892 12396 5058 12420
rect 2980 11720 3000 11780
rect 3120 11720 3324 11780
rect 2980 11700 3324 11720
rect 3770 11680 3840 12380
rect 3620 11640 3840 11680
rect 2360 11540 3540 11622
rect 2180 11328 2320 11420
rect 2360 11414 2560 11540
rect 2960 11480 3140 11502
rect 2960 11400 3000 11480
rect 3080 11400 3140 11480
rect 2348 11328 2562 11360
rect 2180 11280 2562 11328
rect 2960 11280 3140 11400
rect 3440 11420 3540 11540
rect 3620 11520 3660 11640
rect 3718 11520 3840 11640
rect 3620 11480 3840 11520
rect 3440 11340 3616 11420
rect 2180 11240 2740 11280
rect 2180 11182 2560 11240
rect 2700 11182 2740 11240
rect 2960 11220 3500 11280
rect 2180 11152 2740 11182
rect 760 11040 1740 11130
rect 760 10960 1180 11040
rect 1320 10960 1740 11040
rect 760 10880 1740 10960
rect 2180 10880 2354 11152
rect 3420 11102 3500 11220
rect 2398 11048 3500 11102
rect 560 10502 714 10880
rect 1780 10832 2354 10880
rect 1780 10828 2662 10832
rect 2920 10828 3230 10832
rect 1780 10784 3378 10828
rect 1780 10762 3376 10784
rect 1780 10676 3372 10762
rect 750 10602 1744 10674
rect 1920 10670 3372 10676
rect 1920 10660 2662 10670
rect 560 10336 760 10502
rect -2560 9780 -1360 9860
rect -1302 9780 -1120 9860
rect -2560 9680 -1120 9780
rect -902 9760 300 9860
rect -2420 9640 -1120 9680
rect -980 9700 -300 9760
rect -160 9700 60 9760
rect -980 9640 60 9700
rect -2566 8918 -2460 9640
rect 180 9454 242 9580
rect 192 9380 242 9454
rect 188 9360 480 9380
rect 180 9200 480 9360
rect 180 9196 242 9200
rect 192 9100 242 9196
rect 180 8940 242 9100
rect -2566 8756 -2470 8918
rect -1470 8908 120 8912
rect -2424 8792 120 8908
rect -2152 8780 120 8792
rect -938 8778 120 8780
rect -2566 8600 -2180 8756
rect 634 8740 760 10336
rect 1440 10300 1738 10602
rect 1920 10598 2560 10660
rect 1920 10512 2354 10598
rect 1920 10460 2352 10512
rect 3420 10454 3500 11048
rect 3544 10780 3616 11340
rect 3770 11150 3840 11480
rect 3720 11020 3924 11042
rect 3720 10960 3740 11020
rect 3900 10960 3924 11020
rect 4020 11040 5060 11142
rect 4020 10980 4516 11040
rect 4620 10980 5060 11040
rect 4020 10960 5060 10980
rect 3720 10820 3924 10960
rect 3740 10788 3924 10820
rect 3544 10580 3700 10780
rect 3730 10550 3920 10582
rect 2400 10400 3500 10454
rect 3720 10500 3920 10550
rect 3720 10440 3760 10500
rect 3860 10440 3920 10500
rect 3720 10432 3920 10440
rect 3420 10302 3500 10400
rect 3238 10300 3500 10302
rect 3700 10300 3902 10400
rect 1440 10160 3500 10300
rect 158 8520 802 8740
rect 160 7758 200 8520
rect 3238 7740 3500 10160
rect 5260 9858 5320 12440
rect 4020 9820 5322 9858
rect 4020 9720 4040 9820
rect 4180 9720 5322 9820
rect 4020 9682 5322 9720
rect -820 7730 130 7740
rect 240 7730 3940 7740
rect -820 7720 3940 7730
rect -860 7620 3940 7720
rect 4458 5640 5122 5662
rect 4458 5462 4778 5640
rect 5098 5462 5122 5640
rect 4458 5372 5122 5462
rect 5260 5400 5320 9682
rect 5354 5372 6564 5404
rect 4458 5300 6564 5372
rect 4458 5298 5122 5300
<< via1 >>
rect -1200 11940 -1080 12040
rect 460 11940 580 12040
rect 3000 11720 3120 11780
rect 3000 11400 3080 11480
rect 3660 11520 3718 11640
rect 2560 11182 2700 11240
rect 1180 10960 1320 11040
rect -300 9700 -160 9760
rect 3740 10960 3900 11020
rect 4516 10980 4620 11040
rect 3760 10440 3860 10500
rect 4040 9720 4180 9820
rect 4778 5462 5098 5640
<< metal2 >>
rect -1240 12040 600 12080
rect -1240 11940 -1200 12040
rect -1080 11940 460 12040
rect 580 11940 600 12040
rect -1240 11900 600 11940
rect 2980 11780 3140 11802
rect 2980 11720 3000 11780
rect 3120 11720 3140 11780
rect 2980 11480 3140 11720
rect 2980 11400 3000 11480
rect 3080 11400 3140 11480
rect 2980 11380 3140 11400
rect 3640 11640 3740 11680
rect 3640 11520 3660 11640
rect 3718 11520 3740 11640
rect 3640 11260 3740 11520
rect 2540 11240 3740 11260
rect 2540 11182 2560 11240
rect 2700 11182 3740 11240
rect 2540 11160 3740 11182
rect 1160 11040 1340 11060
rect 4480 11040 4660 11080
rect 1160 10960 1180 11040
rect 1320 11020 3922 11040
rect 1320 10960 3740 11020
rect 3900 10960 3922 11020
rect 1160 10940 3922 10960
rect 4480 10980 4516 11040
rect 4620 10980 4660 11040
rect 3740 10500 3872 10506
rect 3740 10440 3760 10500
rect 3860 10440 3872 10500
rect 3740 10400 3872 10440
rect 3700 10380 3902 10400
rect 3700 10320 3760 10380
rect 3860 10320 3902 10380
rect 3700 10300 3902 10320
rect -322 9820 4220 9860
rect -322 9760 4040 9820
rect -322 9700 -300 9760
rect -160 9720 4040 9760
rect 4180 9720 4220 9820
rect -160 9700 4220 9720
rect -322 9682 4220 9700
rect 4480 6000 4660 10980
rect 4480 5740 5182 6000
rect 4480 5682 4760 5740
rect 5100 5682 5182 5740
rect 4480 5640 5182 5682
rect 4480 5570 4778 5640
rect 4754 5462 4778 5570
rect 5098 5462 5182 5640
rect 4754 5438 5182 5462
<< via2 >>
rect 3760 10320 3860 10380
rect 4760 5682 5100 5740
<< metal3 >>
rect 1440 10160 1738 10670
rect 3700 10380 3902 10400
rect 3700 10320 3760 10380
rect 3860 10320 3902 10380
rect 3700 10300 3902 10320
rect 4656 5740 5182 6000
rect 4656 5682 4760 5740
rect 5100 5682 5182 5740
rect 4656 5570 5182 5682
rect 4754 5438 5182 5570
<< metal4 >>
rect 3680 10080 3920 10400
use sky130_fd_pr__cap_mim_m3_1_5JY5WN  XC_c
timestamp 1768734963
transform -1 0 2909 0 -1 7982
box -2370 -2320 2369 2320
use sky130_fd_pr__nfet_01v8_2ZP93L  XM2
timestamp 1768737176
transform 0 -1 -1896 1 0 9276
box -416 -624 416 624
use sky130_fd_pr__pfet_01v8_SZN6ZN  XM4
timestamp 1768735447
transform 0 1 -1922 -1 0 11123
box -1355 -698 1355 664
use sky130_fd_pr__pfet_01v8_B33NDC  XM5
timestamp 1768751538
transform 0 1 2422 -1 0 12351
box -109 -164 109 198
use sky130_fd_pr__nfet_01v8_ND6MQZ  XM8
timestamp 1768749944
transform 0 1 2857 -1 0 10558
box -158 -557 158 557
use sky130_fd_pr__nfet_01v8_73QE7N  XM10
timestamp 1768756364
transform 0 1 -343 -1 0 8245
box -545 -557 545 557
use sky130_fd_pr__pfet_01v8_XL4TZD  XM11
timestamp 1768735973
transform 0 1 1302 -1 0 11758
box -710 -664 710 698
use sky130_fd_pr__nfet_01v8_QG6R6A  XM13
timestamp 1768749944
transform 0 -1 3799 1 0 10686
box -158 -157 158 157
use sky130_fd_pr__pfet_01v8_CYNCWQ  XM14
timestamp 1768736825
transform 0 -1 5926 1 0 8927
box -3605 -698 3605 664
use sky130_fd_pr__nfet_01v8_C8PJZM  XM15
timestamp 1768750829
transform 0 1 4441 -1 0 11768
box -674 -657 674 657
use sky130_fd_pr__nfet_01v8_L4PCGF  sky130_fd_pr__nfet_01v8_L4PCGF_0
timestamp 1768734963
transform 0 1 1248 -1 0 10778
box -158 -588 158 588
use sky130_fd_pr__nfet_01v8_ND6MQZ  sky130_fd_pr__nfet_01v8_ND6MQZ_0
timestamp 1768749944
transform 0 1 2855 -1 0 10938
box -158 -557 158 557
use sky130_fd_pr__nfet_01v8_RYY55T  sky130_fd_pr__nfet_01v8_RYY55T_0
timestamp 1768737176
transform 0 -1 -376 1 0 9276
box -416 -624 416 624
use sky130_fd_pr__pfet_01v8_9WN6ZY  sky130_fd_pr__pfet_01v8_9WN6ZY_0
timestamp 1768735447
transform 0 1 -336 -1 0 11123
box -1355 -664 1355 698
use sky130_fd_pr__pfet_01v8_B33NDC  sky130_fd_pr__pfet_01v8_B33NDC_0
timestamp 1768751538
transform 0 1 2424 -1 0 11869
box -109 -164 109 198
use sky130_fd_pr__pfet_01v8_B33NDC  sky130_fd_pr__pfet_01v8_B33NDC_1
timestamp 1768751538
transform 0 1 2422 -1 0 11387
box -109 -164 109 198
<< labels >>
rlabel metal1 -2566 8600 -2180 8756 0 Vin-
port 9 nsew
rlabel metal1 188 9200 480 9380 0 Vin+
port 10 nsew
rlabel metal1 1920 10460 2352 10880 1 Ptatin
port 11 n
rlabel metal1 3028 11928 3260 12244 1 GND
port 12 n
rlabel metal1 4458 5298 4778 5662 1 Vout
port 13 n
rlabel metal1 -2558 12390 -1358 12800 1 VDD
port 14 n
rlabel space -2558 12390 -1358 12800 1 Vdd
port 15 n
rlabel space -900 12390 300 12800 0 Vsupply
port 16 nsew
<< end >>
