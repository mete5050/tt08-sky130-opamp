magic
tech sky130B
timestamp 1768735072
<< nmos >>
rect -308 -300 -208 300
rect -179 -300 -79 300
rect -50 -300 50 300
rect 79 -300 179 300
rect 208 -300 308 300
<< ndiff >>
rect -337 294 -308 300
rect -337 -294 -331 294
rect -314 -294 -308 294
rect -337 -300 -308 -294
rect -208 294 -179 300
rect -208 -294 -202 294
rect -185 -294 -179 294
rect -208 -300 -179 -294
rect -79 294 -50 300
rect -79 -294 -73 294
rect -56 -294 -50 294
rect -79 -300 -50 -294
rect 50 294 79 300
rect 50 -294 56 294
rect 73 -294 79 294
rect 50 -300 79 -294
rect 179 294 208 300
rect 179 -294 185 294
rect 202 -294 208 294
rect 179 -300 208 -294
rect 308 294 337 300
rect 308 -294 314 294
rect 331 -294 337 294
rect 308 -300 337 -294
<< ndiffc >>
rect -331 -294 -314 294
rect -202 -294 -185 294
rect -73 -294 -56 294
rect 56 -294 73 294
rect 185 -294 202 294
rect 314 -294 331 294
<< poly >>
rect -308 336 -208 344
rect -308 319 -300 336
rect -216 319 -208 336
rect -308 300 -208 319
rect -179 336 -79 344
rect -179 319 -171 336
rect -87 319 -79 336
rect -179 300 -79 319
rect -50 336 50 344
rect -50 319 -42 336
rect 42 319 50 336
rect -50 300 50 319
rect 79 336 179 344
rect 79 319 87 336
rect 171 319 179 336
rect 79 300 179 319
rect 208 336 308 344
rect 208 319 216 336
rect 300 319 308 336
rect 208 300 308 319
rect -308 -319 -208 -300
rect -308 -336 -300 -319
rect -216 -336 -208 -319
rect -308 -344 -208 -336
rect -179 -319 -79 -300
rect -179 -336 -171 -319
rect -87 -336 -79 -319
rect -179 -344 -79 -336
rect -50 -319 50 -300
rect -50 -336 -42 -319
rect 42 -336 50 -319
rect -50 -344 50 -336
rect 79 -319 179 -300
rect 79 -336 87 -319
rect 171 -336 179 -319
rect 79 -344 179 -336
rect 208 -319 308 -300
rect 208 -336 216 -319
rect 300 -336 308 -319
rect 208 -344 308 -336
<< polycont >>
rect -300 319 -216 336
rect -171 319 -87 336
rect -42 319 42 336
rect 87 319 171 336
rect 216 319 300 336
rect -300 -336 -216 -319
rect -171 -336 -87 -319
rect -42 -336 42 -319
rect 87 -336 171 -319
rect 216 -336 300 -319
<< locali >>
rect -308 319 -300 336
rect -216 319 -208 336
rect -179 319 -171 336
rect -87 319 -79 336
rect -50 319 -42 336
rect 42 319 50 336
rect 79 319 87 336
rect 171 319 179 336
rect 208 319 216 336
rect 300 319 308 336
rect -331 294 -314 302
rect -331 -302 -314 -294
rect -202 294 -185 302
rect -202 -302 -185 -294
rect -73 294 -56 302
rect -73 -302 -56 -294
rect 56 294 73 302
rect 56 -302 73 -294
rect 185 294 202 302
rect 185 -302 202 -294
rect 314 294 331 302
rect 314 -302 331 -294
rect -308 -336 -300 -319
rect -216 -336 -208 -319
rect -179 -336 -171 -319
rect -87 -336 -79 -319
rect -50 -336 -42 -319
rect 42 -336 50 -319
rect 79 -336 87 -319
rect 171 -336 179 -319
rect 208 -336 216 -319
rect 300 -336 308 -319
<< viali >>
rect -300 319 -216 336
rect -171 319 -87 336
rect -42 319 42 336
rect 87 319 171 336
rect 216 319 300 336
rect -331 -294 -314 294
rect -202 -294 -185 294
rect -73 -294 -56 294
rect 56 -294 73 294
rect 185 -294 202 294
rect 314 -294 331 294
rect -300 -336 -216 -319
rect -171 -336 -87 -319
rect -42 -336 42 -319
rect 87 -336 171 -319
rect 216 -336 300 -319
<< metal1 >>
rect -306 336 -210 339
rect -306 319 -300 336
rect -216 319 -210 336
rect -306 316 -210 319
rect -177 336 -81 339
rect -177 319 -171 336
rect -87 319 -81 336
rect -177 316 -81 319
rect -48 336 48 339
rect -48 319 -42 336
rect 42 319 48 336
rect -48 316 48 319
rect 81 336 177 339
rect 81 319 87 336
rect 171 319 177 336
rect 81 316 177 319
rect 210 336 306 339
rect 210 319 216 336
rect 300 319 306 336
rect 210 316 306 319
rect -334 294 -311 300
rect -334 -294 -331 294
rect -314 -294 -311 294
rect -334 -300 -311 -294
rect -205 294 -182 300
rect -205 -294 -202 294
rect -185 -294 -182 294
rect -205 -300 -182 -294
rect -76 294 -53 300
rect -76 -294 -73 294
rect -56 -294 -53 294
rect -76 -300 -53 -294
rect 53 294 76 300
rect 53 -294 56 294
rect 73 -294 76 294
rect 53 -300 76 -294
rect 182 294 205 300
rect 182 -294 185 294
rect 202 -294 205 294
rect 182 -300 205 -294
rect 311 294 334 300
rect 311 -294 314 294
rect 331 -294 334 294
rect 311 -300 334 -294
rect -306 -319 -210 -316
rect -306 -336 -300 -319
rect -216 -336 -210 -319
rect -306 -339 -210 -336
rect -177 -319 -81 -316
rect -177 -336 -171 -319
rect -87 -336 -81 -319
rect -177 -339 -81 -336
rect -48 -319 48 -316
rect -48 -336 -42 -319
rect 42 -336 48 -319
rect -48 -339 48 -336
rect 81 -319 177 -316
rect 81 -336 87 -319
rect 171 -336 177 -319
rect 81 -339 177 -336
rect 210 -319 306 -316
rect 210 -336 216 -319
rect 300 -336 306 -319
rect 210 -339 306 -336
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
