magic
tech sky130B
magscale 1 2
timestamp 1768734963
<< nmos >>
rect -358 -567 -158 567
rect -100 -567 100 567
rect 158 -567 358 567
<< ndiff >>
rect -416 555 -358 567
rect -416 -555 -404 555
rect -370 -555 -358 555
rect -416 -567 -358 -555
rect -158 555 -100 567
rect -158 -555 -146 555
rect -112 -555 -100 555
rect -158 -567 -100 -555
rect 100 555 158 567
rect 100 -555 112 555
rect 146 -555 158 555
rect 100 -567 158 -555
rect 358 555 416 567
rect 358 -555 370 555
rect 404 -555 416 555
rect 358 -567 416 -555
<< ndiffc >>
rect -404 -555 -370 555
rect -146 -555 -112 555
rect 112 -555 146 555
rect 370 -555 404 555
<< poly >>
rect -358 639 -158 655
rect -358 605 -342 639
rect -174 605 -158 639
rect -358 567 -158 605
rect -100 639 100 655
rect -100 605 -84 639
rect 84 605 100 639
rect -100 567 100 605
rect 158 639 358 655
rect 158 605 174 639
rect 342 605 358 639
rect 158 567 358 605
rect -358 -605 -158 -567
rect -358 -639 -342 -605
rect -174 -639 -158 -605
rect -358 -655 -158 -639
rect -100 -605 100 -567
rect -100 -639 -84 -605
rect 84 -639 100 -605
rect -100 -655 100 -639
rect 158 -605 358 -567
rect 158 -639 174 -605
rect 342 -639 358 -605
rect 158 -655 358 -639
<< polycont >>
rect -342 605 -174 639
rect -84 605 84 639
rect 174 605 342 639
rect -342 -639 -174 -605
rect -84 -639 84 -605
rect 174 -639 342 -605
<< locali >>
rect -358 605 -342 639
rect -174 605 -158 639
rect -100 605 -84 639
rect 84 605 100 639
rect 158 605 174 639
rect 342 605 358 639
rect -404 555 -370 571
rect -404 -571 -370 -555
rect -146 555 -112 571
rect -146 -571 -112 -555
rect 112 555 146 571
rect 112 -571 146 -555
rect 370 555 404 571
rect 370 -571 404 -555
rect -358 -639 -342 -605
rect -174 -639 -158 -605
rect -100 -639 -84 -605
rect 84 -639 100 -605
rect 158 -639 174 -605
rect 342 -639 358 -605
<< viali >>
rect -342 605 -174 639
rect -84 605 84 639
rect 174 605 342 639
rect -404 -555 -370 555
rect -146 -555 -112 555
rect 112 -555 146 555
rect 370 -555 404 555
rect -342 -639 -174 -605
rect -84 -639 84 -605
rect 174 -639 342 -605
<< metal1 >>
rect -354 639 -162 645
rect -354 605 -342 639
rect -174 605 -162 639
rect -354 599 -162 605
rect -96 639 96 645
rect -96 605 -84 639
rect 84 605 96 639
rect -96 599 96 605
rect 162 639 354 645
rect 162 605 174 639
rect 342 605 354 639
rect 162 599 354 605
rect -410 555 -364 567
rect -410 -555 -404 555
rect -370 -555 -364 555
rect -410 -567 -364 -555
rect -152 555 -106 567
rect -152 -555 -146 555
rect -112 -555 -106 555
rect -152 -567 -106 -555
rect 106 555 152 567
rect 106 -555 112 555
rect 146 -555 152 555
rect 106 -567 152 -555
rect 364 555 410 567
rect 364 -555 370 555
rect 404 -555 410 555
rect 364 -567 410 -555
rect -354 -605 -162 -599
rect -354 -639 -342 -605
rect -174 -639 -162 -605
rect -354 -645 -162 -639
rect -96 -605 96 -599
rect -96 -639 -84 -605
rect 84 -639 96 -605
rect -96 -645 96 -639
rect 162 -605 354 -599
rect 162 -639 174 -605
rect 342 -639 354 -605
rect 162 -645 354 -639
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.666666666666667 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
